// Verilog netlist produced by program LSE :  version Diamond (64-bit) 3.11.2.446
// Netlist written on Sun Sep 13 15:50:56 2020
//
// Verilog Description of module drone2
//

module drone2 (motor_1_pwm, motor_2_pwm, motor_3_pwm, motor_4_pwm, resetn_imu, 
            resetn_lidar, led_data_out, throttle_pwm, yaw_pwm, roll_pwm, 
            pitch_pwm, aux1_pwm, aux2_pwm, swa_swb_pwm, machxo3_switch_reset_n, 
            force_i2c_stall_input_n, sda_1, sda_2, scl_1, scl_2, sin, 
            rxrdy_n, sout, txrdy_n) /* synthesis syn_module_defined=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(42[8:14])
    output motor_1_pwm;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(44[17:28])
    output motor_2_pwm;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(45[17:28])
    output motor_3_pwm;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(46[17:28])
    output motor_4_pwm;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(47[17:28])
    output resetn_imu;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(48[17:27])
    output resetn_lidar;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(49[17:29])
    output [7:0]led_data_out;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(50[23:35])
    input throttle_pwm;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(52[16:28])
    input yaw_pwm;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(53[16:23])
    input roll_pwm;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(54[16:24])
    input pitch_pwm;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(55[16:25])
    input aux1_pwm;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(56[16:24])
    input aux2_pwm;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(57[16:24])
    input swa_swb_pwm;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(58[16:27])
    input machxo3_switch_reset_n;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(59[16:38])
    input force_i2c_stall_input_n;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(60[16:39])
    inout sda_1 /* synthesis black_box_pad_pin=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(62[16:21])
    inout sda_2 /* synthesis black_box_pad_pin=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(63[16:21])
    inout scl_1 /* synthesis black_box_pad_pin=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(64[16:21])
    inout scl_2 /* synthesis black_box_pad_pin=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(65[16:21])
    input sin;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(68[17:20])
    output rxrdy_n;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(69[17:24])
    output sout;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(70[17:21])
    output txrdy_n;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(71[17:24])
    
    wire sys_clk /* synthesis SET_AS_NETWORK=sys_clk, is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(220[10:17])
    wire us_clk /* synthesis SET_AS_NETWORK=us_clk, is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(221[10:16])
    wire sys_clk_N_413 /* synthesis is_inv_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(82[16:24])
    wire i2c2_scli /* synthesis is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_efb_wb.v(34[10:19])
    wire i2c1_scli /* synthesis is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_efb_wb.v(40[10:19])
    
    wire GND_net, motor_1_pwm_c, motor_2_pwm_c, motor_3_pwm_c, motor_4_pwm_c, 
        n17302, led_data_out_c_5, led_data_out_c_4, led_data_out_c_3, 
        led_data_out_c_2, led_data_out_c_1, machxo3_switch_reset_n_c, 
        sin_c, rxrdy_n_c, sout_c;
    wire [7:0]throttle_val;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(76[9:21])
    wire [7:0]yaw_val;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(77[9:16])
    wire [7:0]swa_swb_val;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(82[9:20])
    
    wire n10;
    wire [15:0]next_VL53L1X_chip_id;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(119[9:29])
    wire [15:0]next_VL53L1X_range_mm;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(120[9:30])
    wire [7:0]next_VL53L1X_firm_rdy;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(124[9:30])
    wire [7:0]next_VL53L1X_data_rdy;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(125[9:30])
    wire [7:0]i2c_top_debug_adj_5395;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(53[22:35])
    wire [7:0]next_i2c_device_driver_return_state;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(128[9:44])
    wire [7:0]next_i2c_device_driver_state;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    wire [15:0]VL53L1X_chip_id;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(154[9:24])
    wire [15:0]VL53L1X_range_mm;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(155[9:25])
    wire [7:0]VL53L1X_firm_rdy;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(160[9:25])
    wire [7:0]VL53L1X_data_rdy;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(161[9:25])
    wire [7:0]i2c_device_driver_return_state;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(164[9:39])
    
    wire next_imu_good, next_imu_data_valid;
    wire [7:0]led_data;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(175[16:24])
    
    wire amc_complete_signal;
    wire [15:0]amc_debug;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(184[18:27])
    
    wire throttle_controller_active, resetn;
    wire [1:0]switch_b;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(232[16:24])
    wire [15:0]z_linear_velocity;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(234[17:34])
    wire [7:0]led_data_out_7__N_1;
    
    wire VCC_net;
    wire [7:0]cal_reg_addr;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(105[14:26])
    wire [7:0]next_data_tx_7__N_1032;
    wire [4:0]next_i2c_state_4__N_1055;
    
    wire n8;
    wire [4:0]next_state_4__N_1567;
    
    wire n51135;
    wire [4:0]state_adj_5409;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(74[31:36])
    
    wire count__auto_time_ms_27__N_1639;
    wire [4:0]next_state_4__N_1656;
    wire [8:0]next_auto_state_8__N_1686;
    
    wire next_state_4__N_1666, count__auto_time_ms_27__N_1647;
    wire [6:0]state_adj_5414;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/throttle_controller.v(51[15:20])
    
    wire n48787, n51202, n51186, n51185, n48813, n48828;
    wire [14:0]next_state_14__N_2466;
    
    wire n50715, n48820;
    wire [7:0]latched_pitch;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/angle_controller.v(84[59:72])
    wire [7:0]latched_roll;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/angle_controller.v(84[74:86])
    
    wire n51159, n52179, n36752, n51201, n52, n49185, n50, n48829, 
        n52390, n52389, n34665, n34690, n34692, n52388, n52205, 
        n34474, n38, n37558, high_counter_9__N_4408;
    wire [9:0]next_state_adj_5498;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(92[17:27])
    wire [9:0]state_adj_5499;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(92[29:34])
    wire [3:0]tx_byte_index;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(96[17:30])
    wire [7:0]tx_word_index;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(97[17:30])
    
    wire txrdy_n_c_7, n48722, n49177, n38_adj_5379, n1406;
    wire [15:0]next_dat_i_15__N_4452;
    
    wire state_2__N_199_c_1, n39759, n43309, state_2__N_199_c_1_adj_5380, 
        us_clk_enable_103, state_2__N_199_c_1_adj_5381, n67, n52095, 
        n52092, n43386, state_2__N_199_c_1_adj_5383, wd_event_active, 
        n52359, us_clk_enable_61, byte_rd_left_5__N_1255, n43303, n43302, 
        n27995, n37479, n51044, n41683, n41688, n44, n43271, n33315, 
        n43225, n43221, n43217, n64, n25, n17, n23, n52342, 
        n52341, n49522, n53885;
    wire [2:0]next_state_2__N_4443;
    
    wire i2c2_sdaoen, i2c2_sdao, i2c2_scloen, i2c2_sclo, i2c2_sdai, 
        i2c1_sdaoen, i2c1_sdao, i2c1_scloen, i2c1_sclo, i2c1_sdai, 
        state_2__N_84_c_1, n27, n52142, n123, n27391, n52328, n8774, 
        n36649, n52319, n52318, resetn_derived_2, n52168, n52140, 
        n52306, n4, n50674, n50881, n53884, n15182, n37731, n30695, 
        n52566, n52214, n52213, n51335, n44797, n43332, n52267, 
        n51041, n27734, n52457, n52456, n52441, n51273, n52169, 
        n51272, n51271, n46653, n52429, n48081, n52255;
    
    VHI i2 (.Z(VCC_net));
    FD1S3AX VL53L1X_firm_rdy_i0 (.D(next_VL53L1X_firm_rdy[0]), .CK(sys_clk), 
            .Q(VL53L1X_firm_rdy[0]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_firm_rdy_i0.GSR = "ENABLED";
    FD1S3AX VL53L1X_data_rdy_i0 (.D(next_i2c_state_4__N_1055[1]), .CK(sys_clk), 
            .Q(VL53L1X_data_rdy[0]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_data_rdy_i0.GSR = "ENABLED";
    FD1S3AX led_data_i1 (.D(next_i2c_device_driver_state[0]), .CK(sys_clk), 
            .Q(led_data[0]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam led_data_i1.GSR = "ENABLED";
    FD1S3AX imu_data_valid_78 (.D(next_imu_data_valid), .CK(sys_clk), .Q(next_state_4__N_1567[2]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam imu_data_valid_78.GSR = "ENABLED";
    FD1S3AX imu_good_79 (.D(next_imu_good), .CK(sys_clk), .Q(next_state_14__N_2466[1]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam imu_good_79.GSR = "ENABLED";
    FD1S3AX i2c_device_driver_return_state_i1 (.D(next_i2c_device_driver_return_state[0]), 
            .CK(sys_clk), .Q(i2c_device_driver_return_state[0]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam i2c_device_driver_return_state_i1.GSR = "ENABLED";
    FD1S3AY led_data_out_i1 (.D(led_data_out_7__N_1[1]), .CK(sys_clk), .Q(led_data_out_c_1));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(670[14] 672[12])
    defparam led_data_out_i1.GSR = "ENABLED";
    FD1S3AX resetn_48 (.D(machxo3_switch_reset_n_c), .CK(sys_clk), .Q(resetn));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(567[11] 570[8])
    defparam resetn_48.GSR = "DISABLED";
    OSCH OSCH_inst (.STDBY(GND_net), .OSC(sys_clk)) /* synthesis syn_instantiated=1 */ ;
    defparam OSCH_inst.NOM_FREQ = "38.00";
    OB sout_pad (.I(sout_c), .O(sout));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(70[17:21])
    OB led_data_out_pad_4 (.I(led_data_out_c_4), .O(led_data_out[4]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(50[23:35])
    OB led_data_out_pad_5 (.I(led_data_out_c_5), .O(led_data_out[5]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(50[23:35])
    LUT4 i2c_top_debug_0__bdd_4_lut_40900_4_lut (.A(i2c_top_debug_adj_5395[0]), 
         .B(i2c_top_debug_adj_5395[3]), .C(i2c_top_debug_adj_5395[1]), .D(i2c_top_debug_adj_5395[4]), 
         .Z(n52140)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A ((C+(D))+!B))) */ ;
    defparam i2c_top_debug_0__bdd_4_lut_40900_4_lut.init = 16'h2004;
    OB led_data_out_pad_6 (.I(n17302), .O(led_data_out[6]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(50[23:35])
    ROM256X1A mux_833_Mux_7 (.AD0(cal_reg_addr[0]), .AD1(cal_reg_addr[1]), 
            .AD2(cal_reg_addr[2]), .AD3(cal_reg_addr[3]), .AD4(cal_reg_addr[4]), 
            .AD5(cal_reg_addr[5]), .AD6(cal_reg_addr[6]), .AD7(cal_reg_addr[7]), 
            .DO0(next_data_tx_7__N_1032[7])) /* synthesis initstate=0x0000000000000000000000000000000380008284811000004000000000000000 */ ;
    defparam mux_833_Mux_7.initval = 256'h0000000000000000000000000000000380008284811000004000000000000000;
    ROM256X1A mux_833_Mux_5 (.AD0(cal_reg_addr[0]), .AD1(cal_reg_addr[1]), 
            .AD2(cal_reg_addr[2]), .AD3(cal_reg_addr[3]), .AD4(cal_reg_addr[4]), 
            .AD5(cal_reg_addr[5]), .AD6(cal_reg_addr[6]), .AD7(cal_reg_addr[7]), 
            .DO0(next_data_tx_7__N_1032[5])) /* synthesis initstate=0x0000000000000000000000000000000100000224018010404000000000000000 */ ;
    defparam mux_833_Mux_5.initval = 256'h0000000000000000000000000000000100000224018010404000000000000000;
    ROM256X1A mux_833_Mux_3 (.AD0(cal_reg_addr[0]), .AD1(cal_reg_addr[1]), 
            .AD2(cal_reg_addr[2]), .AD3(cal_reg_addr[3]), .AD4(cal_reg_addr[4]), 
            .AD5(cal_reg_addr[5]), .AD6(cal_reg_addr[6]), .AD7(cal_reg_addr[7]), 
            .DO0(next_data_tx_7__N_1032[3])) /* synthesis initstate=0x000000000000000000000000000000030F00C329899008814050000000000000 */ ;
    defparam mux_833_Mux_3.initval = 256'h000000000000000000000000000000030F00C329899008814050000000000000;
    VLO i1 (.Z(GND_net));
    LUT4 i1_3_lut_4_lut (.A(VL53L1X_chip_id[11]), .B(VL53L1X_chip_id[8]), 
         .C(VL53L1X_chip_id[9]), .D(VL53L1X_chip_id[10]), .Z(n52)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam i1_3_lut_4_lut.init = 16'hfd00;
    ROM256X1A mux_833_Mux_0 (.AD0(cal_reg_addr[0]), .AD1(cal_reg_addr[1]), 
            .AD2(cal_reg_addr[2]), .AD3(cal_reg_addr[3]), .AD4(cal_reg_addr[4]), 
            .AD5(cal_reg_addr[5]), .AD6(cal_reg_addr[6]), .AD7(cal_reg_addr[7]), 
            .DO0(next_data_tx_7__N_1032[0])) /* synthesis initstate=0x0000000000000000000000000000006B8380C01FC30090814301C00000000000 */ ;
    defparam mux_833_Mux_0.initval = 256'h0000000000000000000000000000006B8380C01FC30090814301C00000000000;
    GSR GSR_INST (.GSR(resetn));
    BB BB2_sda (.I(i2c2_sdao), .T(i2c2_sdaoen), .B(sda_2), .O(i2c2_sdai)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=8, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=99, LSE_RLINE=115 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_efb_wb.v(46[8:77])
    BB BB2_scl (.I(i2c2_sclo), .T(i2c2_scloen), .B(scl_2), .O(i2c2_scli)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=8, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=99, LSE_RLINE=115 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_efb_wb.v(48[8:77])
    BB BB1_sda (.I(i2c1_sdao), .T(i2c1_sdaoen), .B(sda_1), .O(i2c1_sdai)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=8, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=99, LSE_RLINE=115 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_efb_wb.v(50[8:77])
    BB BB1_scl (.I(i2c1_sclo), .T(i2c1_scloen), .B(scl_1), .O(i2c1_scli)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=8, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=99, LSE_RLINE=115 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_efb_wb.v(52[8:77])
    OB rxrdy_n_pad (.I(rxrdy_n_c), .O(rxrdy_n));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(69[17:24])
    OB led_data_out_pad_7 (.I(VCC_net), .O(led_data_out[7]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(50[23:35])
    throttle_controller TC (.\state[0] (state_adj_5414[0]), .us_clk(us_clk), 
            .resetn_derived_2(resetn_derived_2), .state({state_adj_5409}), 
            .throttle_controller_active(throttle_controller_active), .resetn(resetn), 
            .n49522(n49522), .\state[2]_adj_6 (state_adj_5414[2]), .\next_state_14__N_2466[1] (next_state_14__N_2466[1]), 
            .n48787(n48787), .n4(n4), .n52214(n52214), .n8(n8), .n30695(n30695), 
            .n8773({n8774}), .n67(n67), .amc_complete_signal(amc_complete_signal), 
            .n37558(n37558), .n39759(n39759), .n52213(n52213), .next_state_4__N_1666(next_state_4__N_1666), 
            .n52566(n52566), .n38(n38_adj_5379)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(377[26] 389[25])
    ROM256X1A mux_833_Mux_2 (.AD0(cal_reg_addr[0]), .AD1(cal_reg_addr[1]), 
            .AD2(cal_reg_addr[2]), .AD3(cal_reg_addr[3]), .AD4(cal_reg_addr[4]), 
            .AD5(cal_reg_addr[5]), .AD6(cal_reg_addr[6]), .AD7(cal_reg_addr[7]), 
            .DO0(next_data_tx_7__N_1032[2])) /* synthesis initstate=0x000000000000000000000000000000018F004009010080014000000000000000 */ ;
    defparam mux_833_Mux_2.initval = 256'h000000000000000000000000000000018F004009010080014000000000000000;
    ROM256X1A mux_833_Mux_1 (.AD0(cal_reg_addr[0]), .AD1(cal_reg_addr[1]), 
            .AD2(cal_reg_addr[2]), .AD3(cal_reg_addr[3]), .AD4(cal_reg_addr[4]), 
            .AD5(cal_reg_addr[5]), .AD6(cal_reg_addr[6]), .AD7(cal_reg_addr[7]), 
            .DO0(next_data_tx_7__N_1032[1])) /* synthesis initstate=0x00000000000000000000000000000043CD00400181000C81400A000000000000 */ ;
    defparam mux_833_Mux_1.initval = 256'h00000000000000000000000000000043CD00400181000C81400A000000000000;
    LUT4 i32806_3_lut_4_lut (.A(i2c_device_driver_return_state[0]), .B(i2c_device_driver_return_state[3]), 
         .C(i2c_device_driver_return_state[1]), .D(i2c_device_driver_return_state[2]), 
         .Z(n43386)) /* synthesis lut_function=(A (C)+!A !(B (C+!(D))+!B !(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam i32806_3_lut_4_lut.init = 16'hb4b0;
    PFUMX i16868 (.BLUT(n48722), .ALUT(n48829), .C0(i2c_top_debug_adj_5395[4]), 
          .Z(n27391));
    LUT4 led_data_6__I_0_i2_1_lut (.A(led_data[0]), .Z(led_data_out_7__N_1[1])) /* synthesis lut_function=(!(A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(671[29:43])
    defparam led_data_6__I_0_i2_1_lut.init = 16'h5555;
    IB sin_pad (.I(sin), .O(sin_c));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(68[17:20])
    IB machxo3_switch_reset_n_pad (.I(machxo3_switch_reset_n), .O(machxo3_switch_reset_n_c));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(59[16:38])
    IB state_2__N_199_pad_1 (.I(swa_swb_pwm), .O(state_2__N_199_c_1_adj_5383));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(58[16:27])
    IB state_2__N_199_pad_1__adj_517 (.I(pitch_pwm), .O(state_2__N_199_c_1_adj_5381));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(55[16:25])
    IB state_2__N_199_pad_1__adj_518 (.I(roll_pwm), .O(state_2__N_199_c_1_adj_5380));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(54[16:24])
    IB state_2__N_199_pad_1__adj_519 (.I(yaw_pwm), .O(state_2__N_199_c_1));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(53[16:23])
    IB state_2__N_84_pad_1 (.I(throttle_pwm), .O(state_2__N_84_c_1));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(52[16:28])
    LUT4 led_data_6__I_0_i5_1_lut_rep_383 (.A(led_data[3]), .Z(n52319)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(671[29:43])
    defparam led_data_6__I_0_i5_1_lut_rep_383.init = 16'h5555;
    LUT4 n42194_bdd_3_lut_40372_4_lut (.A(VL53L1X_range_mm[8]), .B(VL53L1X_range_mm[11]), 
         .C(VL53L1X_range_mm[10]), .D(VL53L1X_range_mm[9]), .Z(n51135)) /* synthesis lut_function=(A (C)+!A (B (C (D))+!B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam n42194_bdd_3_lut_40372_4_lut.init = 16'hf0b0;
    LUT4 n42194_bdd_3_lut_4_lut (.A(VL53L1X_range_mm[8]), .B(VL53L1X_range_mm[11]), 
         .C(VL53L1X_range_mm[9]), .D(VL53L1X_range_mm[10]), .Z(n51335)) /* synthesis lut_function=(A (C)+!A !(B (C+!(D))+!B !(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam n42194_bdd_3_lut_4_lut.init = 16'hb4b0;
    LUT4 i38727_4_lut (.A(throttle_controller_active), .B(n8774), .C(n39759), 
         .D(n67), .Z(n49522)) /* synthesis lut_function=(A (B+!(C+(D)))+!A (B (C+(D)))) */ ;
    defparam i38727_4_lut.init = 16'hccca;
    LUT4 i1_2_lut_rep_331_2_lut (.A(led_data[3]), .B(led_data[1]), .Z(n52267)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(671[29:43])
    defparam i1_2_lut_rep_331_2_lut.init = 16'hdddd;
    LUT4 i1_2_lut_rep_452 (.A(VL53L1X_range_mm[0]), .B(VL53L1X_range_mm[3]), 
         .Z(n52388)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam i1_2_lut_rep_452.init = 16'hbbbb;
    LUT4 i1_3_lut_4_lut_adj_520 (.A(VL53L1X_range_mm[0]), .B(VL53L1X_range_mm[3]), 
         .C(VL53L1X_range_mm[2]), .D(VL53L1X_range_mm[1]), .Z(n25)) /* synthesis lut_function=(A (C)+!A (B (C (D))+!B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam i1_3_lut_4_lut_adj_520.init = 16'hf0b0;
    LUT4 i1_2_lut_rep_453 (.A(VL53L1X_data_rdy[3]), .B(VL53L1X_data_rdy[0]), 
         .Z(n52389)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam i1_2_lut_rep_453.init = 16'hdddd;
    LUT4 i1_3_lut_4_lut_adj_521 (.A(VL53L1X_data_rdy[3]), .B(VL53L1X_data_rdy[0]), 
         .C(VL53L1X_data_rdy[1]), .D(VL53L1X_data_rdy[2]), .Z(n38)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam i1_3_lut_4_lut_adj_521.init = 16'hfd00;
    LUT4 i1_2_lut_rep_454 (.A(VL53L1X_range_mm[4]), .B(VL53L1X_range_mm[7]), 
         .Z(n52390)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam i1_2_lut_rep_454.init = 16'hbbbb;
    LUT4 i7009_2_lut (.A(next_state_2__N_4443[0]), .B(high_counter_9__N_4408), 
         .Z(us_clk_enable_61)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i7009_2_lut.init = 16'hdddd;
    OB resetn_lidar_pad (.I(n52205), .O(resetn_lidar));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(49[17:29])
    OB resetn_imu_pad (.I(n52205), .O(resetn_imu));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(48[17:27])
    OB motor_4_pwm_pad (.I(motor_4_pwm_c), .O(motor_4_pwm));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(47[17:28])
    OB motor_3_pwm_pad (.I(motor_3_pwm_c), .O(motor_3_pwm));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(46[17:28])
    FD1S3AX VL53L1X_chip_id_i0 (.D(next_VL53L1X_chip_id[0]), .CK(sys_clk), 
            .Q(VL53L1X_chip_id[0]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_chip_id_i0.GSR = "ENABLED";
    TSALL TSALL_INST (.TSALL(GND_net));
    LUT4 i1_2_lut_3_lut (.A(VL53L1X_range_mm[2]), .B(VL53L1X_range_mm[1]), 
         .C(VL53L1X_range_mm[3]), .Z(n23)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(155[9:25])
    defparam i1_2_lut_3_lut.init = 16'he0e0;
    LUT4 i14_3_lut_4_lut (.A(VL53L1X_range_mm[2]), .B(VL53L1X_range_mm[1]), 
         .C(VL53L1X_range_mm[3]), .D(VL53L1X_range_mm[0]), .Z(n43225)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B !(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(155[9:25])
    defparam i14_3_lut_4_lut.init = 16'h1fe0;
    LUT4 i1_2_lut_3_lut_adj_522 (.A(VL53L1X_range_mm[6]), .B(VL53L1X_range_mm[5]), 
         .C(VL53L1X_range_mm[7]), .Z(n17)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(155[9:25])
    defparam i1_2_lut_3_lut_adj_522.init = 16'he0e0;
    OB motor_2_pwm_pad (.I(motor_2_pwm_c), .O(motor_2_pwm));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(45[17:28])
    OB motor_1_pwm_pad (.I(motor_1_pwm_c), .O(motor_1_pwm));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(44[17:28])
    LUT4 i11_3_lut_4_lut (.A(VL53L1X_range_mm[6]), .B(VL53L1X_range_mm[5]), 
         .C(VL53L1X_range_mm[7]), .D(VL53L1X_range_mm[4]), .Z(n43221)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B !(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(155[9:25])
    defparam i11_3_lut_4_lut.init = 16'h1fe0;
    PFUMX i32633 (.BLUT(n17), .ALUT(n23), .C0(tx_byte_index[0]), .Z(n43217));
    PUR PUR_INST (.PUR(VCC_net));
    defparam PUR_INST.RST_PULSE = 1;
    LUT4 i1_2_lut (.A(VL53L1X_data_rdy[7]), .B(VL53L1X_data_rdy[4]), .Z(n34474)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam i1_2_lut.init = 16'hdddd;
    FD1S3AX led_data_out_i6 (.D(n53885), .CK(sys_clk), .Q(n17302));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(670[14] 672[12])
    defparam led_data_out_i6.GSR = "ENABLED";
    FD1S3AY led_data_out_i5 (.D(led_data_out_7__N_1[5]), .CK(sys_clk), .Q(led_data_out_c_5));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(670[14] 672[12])
    defparam led_data_out_i5.GSR = "ENABLED";
    FD1S3AX led_data_out_i4 (.D(n52319), .CK(sys_clk), .Q(led_data_out_c_4));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(670[14] 672[12])
    defparam led_data_out_i4.GSR = "ENABLED";
    FD1S3AY led_data_out_i3 (.D(led_data_out_7__N_1[3]), .CK(sys_clk), .Q(led_data_out_c_3));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(670[14] 672[12])
    defparam led_data_out_i3.GSR = "ENABLED";
    FD1S3AX led_data_out_i2 (.D(led_data_out_7__N_1[2]), .CK(sys_clk), .Q(led_data_out_c_2));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(670[14] 672[12])
    defparam led_data_out_i2.GSR = "ENABLED";
    FD1S3AX i2c_device_driver_return_state_i5 (.D(next_i2c_device_driver_return_state[4]), 
            .CK(sys_clk), .Q(i2c_device_driver_return_state[4]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam i2c_device_driver_return_state_i5.GSR = "ENABLED";
    FD1S3AX i2c_device_driver_return_state_i4 (.D(next_i2c_device_driver_return_state[3]), 
            .CK(sys_clk), .Q(i2c_device_driver_return_state[3]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam i2c_device_driver_return_state_i4.GSR = "ENABLED";
    FD1S3AX i2c_device_driver_return_state_i3 (.D(next_i2c_device_driver_return_state[2]), 
            .CK(sys_clk), .Q(i2c_device_driver_return_state[2]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam i2c_device_driver_return_state_i3.GSR = "ENABLED";
    FD1S3AX i2c_device_driver_return_state_i2 (.D(next_i2c_device_driver_return_state[1]), 
            .CK(sys_clk), .Q(i2c_device_driver_return_state[1]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam i2c_device_driver_return_state_i2.GSR = "ENABLED";
    FD1S3AX led_data_i5 (.D(next_i2c_device_driver_state[4]), .CK(sys_clk), 
            .Q(led_data[4]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam led_data_i5.GSR = "ENABLED";
    FD1S3AX led_data_i4 (.D(next_i2c_device_driver_state[3]), .CK(sys_clk), 
            .Q(led_data[3]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam led_data_i4.GSR = "ENABLED";
    FD1S3AX led_data_i3 (.D(next_i2c_device_driver_state[2]), .CK(sys_clk), 
            .Q(led_data[2]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam led_data_i3.GSR = "ENABLED";
    FD1S3AX led_data_i2 (.D(next_i2c_device_driver_state[1]), .CK(sys_clk), 
            .Q(led_data[1]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam led_data_i2.GSR = "ENABLED";
    FD1S3AX VL53L1X_data_rdy_i7 (.D(next_VL53L1X_data_rdy[7]), .CK(sys_clk), 
            .Q(VL53L1X_data_rdy[7]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_data_rdy_i7.GSR = "ENABLED";
    FD1S3AX VL53L1X_data_rdy_i6 (.D(next_VL53L1X_data_rdy[6]), .CK(sys_clk), 
            .Q(VL53L1X_data_rdy[6]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_data_rdy_i6.GSR = "ENABLED";
    FD1S3AX VL53L1X_data_rdy_i5 (.D(next_VL53L1X_data_rdy[5]), .CK(sys_clk), 
            .Q(VL53L1X_data_rdy[5]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_data_rdy_i5.GSR = "ENABLED";
    FD1S3AX VL53L1X_data_rdy_i4 (.D(next_VL53L1X_data_rdy[4]), .CK(sys_clk), 
            .Q(VL53L1X_data_rdy[4]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_data_rdy_i4.GSR = "ENABLED";
    FD1S3AX VL53L1X_data_rdy_i3 (.D(next_VL53L1X_data_rdy[3]), .CK(sys_clk), 
            .Q(VL53L1X_data_rdy[3]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_data_rdy_i3.GSR = "ENABLED";
    FD1S3AX VL53L1X_data_rdy_i2 (.D(next_VL53L1X_data_rdy[2]), .CK(sys_clk), 
            .Q(VL53L1X_data_rdy[2]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_data_rdy_i2.GSR = "ENABLED";
    FD1S3AX VL53L1X_data_rdy_i1 (.D(next_VL53L1X_data_rdy[1]), .CK(sys_clk), 
            .Q(VL53L1X_data_rdy[1]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_data_rdy_i1.GSR = "ENABLED";
    FD1S3AX VL53L1X_firm_rdy_i7 (.D(next_VL53L1X_firm_rdy[7]), .CK(sys_clk), 
            .Q(VL53L1X_firm_rdy[7]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_firm_rdy_i7.GSR = "ENABLED";
    FD1S3AX VL53L1X_firm_rdy_i6 (.D(next_VL53L1X_firm_rdy[6]), .CK(sys_clk), 
            .Q(VL53L1X_firm_rdy[6]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_firm_rdy_i6.GSR = "ENABLED";
    FD1S3AX VL53L1X_firm_rdy_i5 (.D(next_VL53L1X_firm_rdy[5]), .CK(sys_clk), 
            .Q(VL53L1X_firm_rdy[5]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_firm_rdy_i5.GSR = "ENABLED";
    FD1S3AX VL53L1X_firm_rdy_i4 (.D(next_VL53L1X_firm_rdy[4]), .CK(sys_clk), 
            .Q(VL53L1X_firm_rdy[4]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_firm_rdy_i4.GSR = "ENABLED";
    FD1S3AX VL53L1X_firm_rdy_i3 (.D(next_VL53L1X_firm_rdy[3]), .CK(sys_clk), 
            .Q(VL53L1X_firm_rdy[3]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_firm_rdy_i3.GSR = "ENABLED";
    FD1S3AX VL53L1X_firm_rdy_i2 (.D(next_VL53L1X_firm_rdy[2]), .CK(sys_clk), 
            .Q(VL53L1X_firm_rdy[2]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_firm_rdy_i2.GSR = "ENABLED";
    FD1S3AX VL53L1X_firm_rdy_i1 (.D(next_VL53L1X_firm_rdy[1]), .CK(sys_clk), 
            .Q(VL53L1X_firm_rdy[1]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_firm_rdy_i1.GSR = "ENABLED";
    FD1S3AX VL53L1X_range_mm_i15 (.D(next_VL53L1X_range_mm[15]), .CK(sys_clk), 
            .Q(VL53L1X_range_mm[15]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_range_mm_i15.GSR = "ENABLED";
    FD1S3AX VL53L1X_range_mm_i14 (.D(next_VL53L1X_range_mm[14]), .CK(sys_clk), 
            .Q(VL53L1X_range_mm[14]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_range_mm_i14.GSR = "ENABLED";
    FD1S3AX VL53L1X_range_mm_i13 (.D(next_VL53L1X_range_mm[13]), .CK(sys_clk), 
            .Q(VL53L1X_range_mm[13]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_range_mm_i13.GSR = "ENABLED";
    FD1S3AX VL53L1X_range_mm_i12 (.D(next_VL53L1X_range_mm[12]), .CK(sys_clk), 
            .Q(VL53L1X_range_mm[12]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_range_mm_i12.GSR = "ENABLED";
    FD1S3AX VL53L1X_range_mm_i11 (.D(next_VL53L1X_range_mm[11]), .CK(sys_clk), 
            .Q(VL53L1X_range_mm[11]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_range_mm_i11.GSR = "ENABLED";
    OB txrdy_n_pad (.I(txrdy_n_c_7), .O(txrdy_n));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(71[17:24])
    FD1S3AX VL53L1X_range_mm_i10 (.D(next_VL53L1X_range_mm[10]), .CK(sys_clk), 
            .Q(VL53L1X_range_mm[10]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_range_mm_i10.GSR = "ENABLED";
    FD1S3AX VL53L1X_range_mm_i9 (.D(next_VL53L1X_range_mm[9]), .CK(sys_clk), 
            .Q(VL53L1X_range_mm[9]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_range_mm_i9.GSR = "ENABLED";
    LUT4 VL53L1X_range_mm_2__bdd_3_lut_40280 (.A(VL53L1X_range_mm[2]), .B(VL53L1X_range_mm[3]), 
         .C(VL53L1X_range_mm[1]), .Z(n51185)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam VL53L1X_range_mm_2__bdd_3_lut_40280.init = 16'h0404;
    LUT4 VL53L1X_range_mm_2__bdd_3_lut (.A(VL53L1X_range_mm[5]), .B(VL53L1X_range_mm[6]), 
         .C(VL53L1X_range_mm[7]), .Z(n51186)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam VL53L1X_range_mm_2__bdd_3_lut.init = 16'h1010;
    FD1S3AX VL53L1X_range_mm_i8 (.D(next_VL53L1X_range_mm[8]), .CK(sys_clk), 
            .Q(VL53L1X_range_mm[8]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_range_mm_i8.GSR = "ENABLED";
    FD1S3AX VL53L1X_range_mm_i7 (.D(next_VL53L1X_range_mm[7]), .CK(sys_clk), 
            .Q(VL53L1X_range_mm[7]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_range_mm_i7.GSR = "ENABLED";
    FD1S3AX VL53L1X_range_mm_i6 (.D(next_VL53L1X_range_mm[6]), .CK(sys_clk), 
            .Q(VL53L1X_range_mm[6]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_range_mm_i6.GSR = "ENABLED";
    FD1S3AX VL53L1X_range_mm_i5 (.D(next_VL53L1X_range_mm[5]), .CK(sys_clk), 
            .Q(VL53L1X_range_mm[5]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_range_mm_i5.GSR = "ENABLED";
    FD1S3AX VL53L1X_range_mm_i4 (.D(next_VL53L1X_range_mm[4]), .CK(sys_clk), 
            .Q(VL53L1X_range_mm[4]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_range_mm_i4.GSR = "ENABLED";
    FD1S3AX VL53L1X_range_mm_i3 (.D(next_VL53L1X_range_mm[3]), .CK(sys_clk), 
            .Q(VL53L1X_range_mm[3]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_range_mm_i3.GSR = "ENABLED";
    FD1S3AX VL53L1X_range_mm_i2 (.D(next_VL53L1X_range_mm[2]), .CK(sys_clk), 
            .Q(VL53L1X_range_mm[2]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_range_mm_i2.GSR = "ENABLED";
    FD1S3AX VL53L1X_range_mm_i1 (.D(next_VL53L1X_range_mm[1]), .CK(sys_clk), 
            .Q(VL53L1X_range_mm[1]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_range_mm_i1.GSR = "ENABLED";
    FD1S3AX VL53L1X_chip_id_i15 (.D(next_VL53L1X_chip_id[15]), .CK(sys_clk), 
            .Q(VL53L1X_chip_id[15]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_chip_id_i15.GSR = "ENABLED";
    FD1S3AX VL53L1X_chip_id_i14 (.D(next_VL53L1X_chip_id[14]), .CK(sys_clk), 
            .Q(VL53L1X_chip_id[14]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_chip_id_i14.GSR = "ENABLED";
    FD1S3AX VL53L1X_chip_id_i13 (.D(next_VL53L1X_chip_id[13]), .CK(sys_clk), 
            .Q(VL53L1X_chip_id[13]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_chip_id_i13.GSR = "ENABLED";
    FD1S3AX VL53L1X_chip_id_i12 (.D(next_VL53L1X_chip_id[12]), .CK(sys_clk), 
            .Q(VL53L1X_chip_id[12]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_chip_id_i12.GSR = "ENABLED";
    FD1S3AX VL53L1X_chip_id_i11 (.D(next_VL53L1X_chip_id[11]), .CK(sys_clk), 
            .Q(VL53L1X_chip_id[11]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_chip_id_i11.GSR = "ENABLED";
    FD1S3AX VL53L1X_chip_id_i10 (.D(next_VL53L1X_chip_id[10]), .CK(sys_clk), 
            .Q(VL53L1X_chip_id[10]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_chip_id_i10.GSR = "ENABLED";
    FD1S3AX VL53L1X_chip_id_i9 (.D(next_VL53L1X_chip_id[9]), .CK(sys_clk), 
            .Q(VL53L1X_chip_id[9]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_chip_id_i9.GSR = "ENABLED";
    FD1S3AX VL53L1X_chip_id_i8 (.D(next_VL53L1X_chip_id[8]), .CK(sys_clk), 
            .Q(VL53L1X_chip_id[8]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_chip_id_i8.GSR = "ENABLED";
    FD1S3AX VL53L1X_chip_id_i7 (.D(next_VL53L1X_chip_id[7]), .CK(sys_clk), 
            .Q(VL53L1X_chip_id[7]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_chip_id_i7.GSR = "ENABLED";
    FD1S3AX VL53L1X_chip_id_i6 (.D(next_VL53L1X_chip_id[6]), .CK(sys_clk), 
            .Q(VL53L1X_chip_id[6]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_chip_id_i6.GSR = "ENABLED";
    FD1S3AX VL53L1X_chip_id_i5 (.D(next_VL53L1X_chip_id[5]), .CK(sys_clk), 
            .Q(VL53L1X_chip_id[5]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_chip_id_i5.GSR = "ENABLED";
    FD1S3AX VL53L1X_chip_id_i4 (.D(next_VL53L1X_chip_id[4]), .CK(sys_clk), 
            .Q(VL53L1X_chip_id[4]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_chip_id_i4.GSR = "ENABLED";
    OB led_data_out_pad_0 (.I(n17302), .O(led_data_out[0]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(50[23:35])
    OB led_data_out_pad_1 (.I(led_data_out_c_1), .O(led_data_out[1]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(50[23:35])
    FD1S3AX VL53L1X_chip_id_i3 (.D(next_VL53L1X_chip_id[3]), .CK(sys_clk), 
            .Q(VL53L1X_chip_id[3]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_chip_id_i3.GSR = "ENABLED";
    OB led_data_out_pad_2 (.I(led_data_out_c_2), .O(led_data_out[2]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(50[23:35])
    FD1S3AX VL53L1X_chip_id_i2 (.D(next_VL53L1X_chip_id[2]), .CK(sys_clk), 
            .Q(VL53L1X_chip_id[2]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_chip_id_i2.GSR = "ENABLED";
    FD1S3AX VL53L1X_chip_id_i1 (.D(next_VL53L1X_chip_id[1]), .CK(sys_clk), 
            .Q(VL53L1X_chip_id[1]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_chip_id_i1.GSR = "ENABLED";
    OB led_data_out_pad_3 (.I(led_data_out_c_3), .O(led_data_out[3]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(50[23:35])
    LUT4 n51186_bdd_4_lut (.A(n51186), .B(n51185), .C(tx_byte_index[0]), 
         .D(tx_byte_index[1]), .Z(n52169)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam n51186_bdd_4_lut.init = 16'hffca;
    LUT4 i2_3_lut (.A(VL53L1X_chip_id[9]), .B(VL53L1X_chip_id[11]), .C(VL53L1X_chip_id[10]), 
         .Z(n49185)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i2_3_lut.init = 16'h0404;
    LUT4 i2_3_lut_adj_523 (.A(VL53L1X_chip_id[14]), .B(VL53L1X_chip_id[13]), 
         .C(VL53L1X_chip_id[15]), .Z(n48828)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i2_3_lut_adj_523.init = 16'h1010;
    LUT4 i1_2_lut_adj_524 (.A(resetn), .B(n67), .Z(n38_adj_5379)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(567[11] 570[8])
    defparam i1_2_lut_adj_524.init = 16'h8888;
    us_clk us_clk_divider (.GND_net(GND_net), .us_clk(us_clk), .sys_clk(sys_clk)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(249[12] 252[25])
    LUT4 i3_4_lut (.A(resetn), .B(n8), .C(state_adj_5414[2]), .D(state_adj_5414[0]), 
         .Z(n30695)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(567[11] 570[8])
    defparam i3_4_lut.init = 16'h0008;
    LUT4 m1_lut (.Z(n53885)) /* synthesis lut_function=1, syn_instantiated=1 */ ;
    defparam m1_lut.init = 16'hffff;
    INV i41687 (.A(sys_clk), .Z(sys_clk_N_413));
    receiver receiver (.state_2__N_199_c_1(state_2__N_199_c_1), .us_clk(us_clk), 
            .GND_net(GND_net), .yaw_val({yaw_val}), .n43271(n43271), .n52456(n52456), 
            .n51041(n51041), .state_2__N_84_c_1(state_2__N_84_c_1), .resetn(resetn), 
            .resetn_derived_2(resetn_derived_2), .\i2c_top_debug[1] (i2c_top_debug_adj_5395[1]), 
            .n52306(n52306), .wd_event_active(wd_event_active), .n52205(n52205), 
            .n44(n44), .n44797(n44797), .n64(n64), .\next_state[0] (next_state_adj_5498[0]), 
            .n33315(n33315), .count__auto_time_ms_27__N_1639(count__auto_time_ms_27__N_1639), 
            .n52318(n52318), .n52142(n52142), .\i2c_top_debug[5] (i2c_top_debug_adj_5395[5]), 
            .byte_rd_left_5__N_1255(byte_rd_left_5__N_1255), .throttle_val({throttle_val}), 
            .n52441(n52441), .n51044(n51044), .n52429(n52429), .swa_swb_val({swa_swb_val}), 
            .state_2__N_199_c_1_adj_2(state_2__N_199_c_1_adj_5383), .state_2__N_199_c_1_adj_3(state_2__N_199_c_1_adj_5380), 
            .\latched_roll[7] (latched_roll[7]), .\latched_roll[6] (latched_roll[6]), 
            .\latched_roll[5] (latched_roll[5]), .\latched_roll[4] (latched_roll[4]), 
            .\latched_roll[2] (latched_roll[2]), .n48820(n48820), .state_2__N_199_c_1_adj_4(state_2__N_199_c_1_adj_5381), 
            .n1406(n1406), .latched_pitch({latched_pitch}), .n52328(n52328), 
            .\tx_byte_index[0] (tx_byte_index[0]), .n52095(n52095), .n27(n27), 
            .\tx_byte_index[1] (tx_byte_index[1]), .\tx_word_index[1] (tx_word_index[1]), 
            .n36649(n36649), .n34665(n34665), .n51272(n51272), .n51271(n51271), 
            .n51273(n51273), .n51202(n51202), .n51159(n51159), .n51201(n51201), 
            .n34692(n34692), .n36752(n36752), .n34690(n34690)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(258[14] 276[25])
    LUT4 m0_lut (.Z(n53884)) /* synthesis lut_function=0, syn_instantiated=1 */ ;
    defparam m0_lut.init = 16'h0000;
    \i2c_device_driver(INIT_INTERVAL=16'b01111101000,POLL_INTERVAL=16'b010100)  I2C_Devices (.sys_clk_N_413(sys_clk_N_413), 
            .sys_clk(sys_clk), .\next_i2c_state_4__N_1055[1] (next_i2c_state_4__N_1055[1]), 
            .\next_i2c_device_driver_state[3] (next_i2c_device_driver_state[3]), 
            .\next_i2c_device_driver_state[2] (next_i2c_device_driver_state[2]), 
            .\next_i2c_device_driver_state[0] (next_i2c_device_driver_state[0]), 
            .\next_i2c_device_driver_state[4] (next_i2c_device_driver_state[4]), 
            .cal_reg_addr({cal_reg_addr}), .resetn(resetn), .next_VL53L1X_firm_rdy({next_VL53L1X_firm_rdy}), 
            .\next_i2c_device_driver_return_state[0] (next_i2c_device_driver_return_state[0]), 
            .n53885(n53885), .next_imu_good(next_imu_good), .\next_i2c_device_driver_return_state[2] (next_i2c_device_driver_return_state[2]), 
            .next_VL53L1X_range_mm({next_VL53L1X_range_mm}), .next_data_tx_7__N_1032({next_data_tx_7__N_1032[7], 
            Open_0, next_data_tx_7__N_1032[5], Open_1, next_data_tx_7__N_1032[3:2], 
            Open_2, next_data_tx_7__N_1032[0]}), .\next_VL53L1X_data_rdy[7] (next_VL53L1X_data_rdy[7]), 
            .next_VL53L1X_chip_id({next_VL53L1X_chip_id}), .\next_VL53L1X_data_rdy[6] (next_VL53L1X_data_rdy[6]), 
            .\i2c_top_debug[1] (i2c_top_debug_adj_5395[1]), .wd_event_active(wd_event_active), 
            .n52306(n52306), .\next_VL53L1X_data_rdy[5] (next_VL53L1X_data_rdy[5]), 
            .\next_VL53L1X_data_rdy[4] (next_VL53L1X_data_rdy[4]), .\next_VL53L1X_data_rdy[3] (next_VL53L1X_data_rdy[3]), 
            .\next_VL53L1X_data_rdy[2] (next_VL53L1X_data_rdy[2]), .\next_VL53L1X_data_rdy[1] (next_VL53L1X_data_rdy[1]), 
            .GND_net(GND_net), .\next_i2c_device_driver_return_state[4] (next_i2c_device_driver_return_state[4]), 
            .\next_i2c_device_driver_return_state[3] (next_i2c_device_driver_return_state[3]), 
            .\next_i2c_device_driver_return_state[1] (next_i2c_device_driver_return_state[1]), 
            .n52205(n52205), .n52318(n52318), .\i2c_top_debug[3] (i2c_top_debug_adj_5395[3]), 
            .\i2c_top_debug[4] (i2c_top_debug_adj_5395[4]), .\next_i2c_device_driver_state[1] (next_i2c_device_driver_state[1]), 
            .throttle_controller_active(throttle_controller_active), .next_imu_data_valid(next_imu_data_valid), 
            .\next_data_tx_7__N_1032[1] (next_data_tx_7__N_1032[1]), .\i2c_top_debug[0] (i2c_top_debug_adj_5395[0]), 
            .\i2c_top_debug[5] (i2c_top_debug_adj_5395[5]), .resetn_derived_2(resetn_derived_2), 
            .byte_rd_left_5__N_1255(byte_rd_left_5__N_1255), .n52142(n52142), 
            .n27391(n27391), .n48722(n48722), .n48829(n48829), .n52140(n52140), 
            .i2c2_sdaoen(i2c2_sdaoen), .i2c2_sdao(i2c2_sdao), .i2c2_scloen(i2c2_scloen), 
            .i2c2_sclo(i2c2_sclo), .i2c2_sdai(i2c2_sdai), .i2c2_scli(i2c2_scli), 
            .i2c1_sdaoen(i2c1_sdaoen), .i2c1_sdao(i2c1_sdao), .i2c1_scloen(i2c1_scloen), 
            .i2c1_sclo(i2c1_sclo), .i2c1_sdai(i2c1_sdai), .i2c1_scli(i2c1_scli), 
            .VCC_net(VCC_net)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(299[9] 349[6])
    LUT4 n38079_bdd_3_lut_40904_4_lut (.A(i2c_device_driver_return_state[1]), 
         .B(i2c_device_driver_return_state[3]), .C(tx_byte_index[0]), .D(i2c_device_driver_return_state[2]), 
         .Z(n52092)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam n38079_bdd_3_lut_40904_4_lut.init = 16'h0040;
    LUT4 i26017_3_lut_4_lut (.A(i2c_device_driver_return_state[1]), .B(i2c_device_driver_return_state[3]), 
         .C(i2c_device_driver_return_state[2]), .D(i2c_device_driver_return_state[0]), 
         .Z(n36649)) /* synthesis lut_function=(A (C)+!A (B (C (D))+!B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam i26017_3_lut_4_lut.init = 16'hf0b0;
    LUT4 led_data_6__I_0_i6_1_lut (.A(led_data[4]), .Z(led_data_out_7__N_1[5])) /* synthesis lut_function=(!(A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(671[29:43])
    defparam led_data_6__I_0_i6_1_lut.init = 16'h5555;
    LUT4 led_data_6__I_0_i4_1_lut (.A(led_data[2]), .Z(led_data_out_7__N_1[3])) /* synthesis lut_function=(!(A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(671[29:43])
    defparam led_data_6__I_0_i4_1_lut.init = 16'h5555;
    LUT4 i2_3_lut_adj_525 (.A(VL53L1X_data_rdy[6]), .B(VL53L1X_data_rdy[5]), 
         .C(VL53L1X_data_rdy[7]), .Z(n48813)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i2_3_lut_adj_525.init = 16'h1010;
    LUT4 i1_2_lut_adj_526 (.A(resetn), .B(n33315), .Z(count__auto_time_ms_27__N_1647)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(567[11] 570[8])
    defparam i1_2_lut_adj_526.init = 16'h8888;
    LUT4 i2_3_lut_adj_527 (.A(VL53L1X_data_rdy[1]), .B(VL53L1X_data_rdy[3]), 
         .C(VL53L1X_data_rdy[2]), .Z(n49177)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i2_3_lut_adj_527.init = 16'h0404;
    LUT4 i1_2_lut_rep_521 (.A(i2c_device_driver_return_state[1]), .B(i2c_device_driver_return_state[2]), 
         .Z(n52457)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(164[9:39])
    defparam i1_2_lut_rep_521.init = 16'heeee;
    LUT4 n18_bdd_3_lut_4_lut (.A(i2c_device_driver_return_state[1]), .B(i2c_device_driver_return_state[2]), 
         .C(i2c_device_driver_return_state[3]), .D(tx_byte_index[0]), .Z(n50881)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(164[9:39])
    defparam n18_bdd_3_lut_4_lut.init = 16'he000;
    LUT4 i1_3_lut_4_lut_adj_528 (.A(VL53L1X_chip_id[12]), .B(VL53L1X_chip_id[15]), 
         .C(VL53L1X_chip_id[13]), .D(VL53L1X_chip_id[14]), .Z(n50)) /* synthesis lut_function=(A (D)+!A (B (C (D))+!B (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam i1_3_lut_4_lut_adj_528.init = 16'hfb00;
    LUT4 tx_byte_index_0__bdd_3_lut_40618_4_lut (.A(VL53L1X_chip_id[11]), 
         .B(VL53L1X_chip_id[8]), .C(VL53L1X_chip_id[10]), .D(VL53L1X_chip_id[9]), 
         .Z(n50674)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A (D)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam tx_byte_index_0__bdd_3_lut_40618_4_lut.init = 16'hdd20;
    z_linear_velocity_comp ZLV (.n53884(n53884), .sys_clk(sys_clk), .\next_state_4__N_1567[2] (next_state_4__N_1567[2]), 
            .\z_linear_velocity[3] (z_linear_velocity[3]), .\z_linear_velocity[1] (z_linear_velocity[1]), 
            .\z_linear_velocity[2] (z_linear_velocity[2]), .n50715(n50715), 
            .\z_linear_velocity[6] (z_linear_velocity[6]), .\z_linear_velocity[5] (z_linear_velocity[5]), 
            .\z_linear_velocity[7] (z_linear_velocity[7]), .\z_linear_velocity[4] (z_linear_velocity[4]), 
            .n43332(n43332), .GND_net(GND_net), .\tx_byte_index[0] (tx_byte_index[0]), 
            .\tx_byte_index[1] (tx_byte_index[1]), .n52168(n52168), .n43302(n43302), 
            .n43303(n43303), .n27734(n27734), .n48081(n48081), .n123(n123), 
            .n52255(n52255), .\next_dat_i_15__N_4452[3] (next_dat_i_15__N_4452[3]), 
            .\next_state_4__N_1656[2] (next_state_4__N_1656[2]), .us_clk_enable_103(us_clk_enable_103), 
            .n46653(n46653), .n52341(n52341), .n37731(n37731), .n52342(n52342), 
            .n15182(n15182), .\state[2] (state_adj_5499[2]), .\state[5] (state_adj_5499[5]), 
            .n43309(n43309), .\z_linear_velocity[10] (z_linear_velocity[10]), 
            .\z_linear_velocity[11] (z_linear_velocity[11]), .\VL53L1X_range_mm[1] (VL53L1X_range_mm[1]), 
            .\VL53L1X_range_mm[2] (VL53L1X_range_mm[2]), .\VL53L1X_range_mm[3] (VL53L1X_range_mm[3]), 
            .\VL53L1X_range_mm[4] (VL53L1X_range_mm[4]), .\VL53L1X_range_mm[5] (VL53L1X_range_mm[5]), 
            .\VL53L1X_range_mm[6] (VL53L1X_range_mm[6]), .\VL53L1X_range_mm[7] (VL53L1X_range_mm[7]), 
            .\VL53L1X_range_mm[8] (VL53L1X_range_mm[8]), .\VL53L1X_range_mm[9] (VL53L1X_range_mm[9]), 
            .\VL53L1X_range_mm[10] (VL53L1X_range_mm[10]), .\VL53L1X_range_mm[11] (VL53L1X_range_mm[11]), 
            .\VL53L1X_range_mm[12] (VL53L1X_range_mm[12]), .\VL53L1X_range_mm[13] (VL53L1X_range_mm[13]), 
            .\VL53L1X_range_mm[14] (VL53L1X_range_mm[14]), .\z_linear_velocity[12] (z_linear_velocity[12]), 
            .\z_linear_velocity[13] (z_linear_velocity[13]), .\z_linear_velocity[14] (z_linear_velocity[14]), 
            .\z_linear_velocity[15] (z_linear_velocity[15]), .\VL53L1X_range_mm[0] (VL53L1X_range_mm[0]), 
            .\z_linear_velocity[8] (z_linear_velocity[8]), .\z_linear_velocity[9] (z_linear_velocity[9])) /* synthesis syn_module_defined=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(352[28] 358[6])
    auto_mode_controller AMC (.state({state_adj_5409}), .resetn_derived_2(resetn_derived_2), 
            .count__auto_time_ms_27__N_1647(count__auto_time_ms_27__N_1647), 
            .n53885(n53885), .us_clk(us_clk), .amc_complete_signal(amc_complete_signal), 
            .\amc_debug[0] (amc_debug[0]), .next_state_4__N_1666(next_state_4__N_1666), 
            .GND_net(GND_net), .\next_state_14__N_2466[1] (next_state_14__N_2466[1]), 
            .\next_state_4__N_1656[2] (next_state_4__N_1656[2]), .n52214(n52214), 
            .n4(n4), .us_clk_enable_103(us_clk_enable_103), .\throttle_val[1] (throttle_val[1]), 
            .switch_b({switch_b}), .\next_auto_state_8__N_1686[7] (next_auto_state_8__N_1686[7]), 
            .\amc_debug[8] (amc_debug[8]), .\amc_debug[7] (amc_debug[7]), 
            .\amc_debug[6] (amc_debug[6]), .\amc_debug[5] (amc_debug[5]), 
            .\amc_debug[4] (amc_debug[4]), .\amc_debug[3] (amc_debug[3]), 
            .\amc_debug[2] (amc_debug[2]), .\amc_debug[1] (amc_debug[1]), 
            .count__auto_time_ms_27__N_1639(count__auto_time_ms_27__N_1639), 
            .n41683(n41683), .n41688(n41688), .n46653(n46653), .\throttle_val[2] (throttle_val[2]), 
            .\throttle_val[3] (throttle_val[3]), .\throttle_val[4] (throttle_val[4]), 
            .\throttle_val[5] (throttle_val[5]), .\throttle_val[6] (throttle_val[6]), 
            .\throttle_val[7] (throttle_val[7]), .n52213(n52213), .n48787(n48787), 
            .n37558(n37558), .n33315(n33315), .n52566(n52566)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(362[26] 375[6])
    flight_mode MODE (.switch_b({switch_b}), .us_clk(us_clk), .\swa_swb_val[7] (swa_swb_val[7]), 
            .\swa_swb_val[4] (swa_swb_val[4]), .\swa_swb_val[5] (swa_swb_val[5]), 
            .\swa_swb_val[3] (swa_swb_val[3]), .\swa_swb_val[6] (swa_swb_val[6]), 
            .\swa_swb_val[2] (swa_swb_val[2]), .n10(n10), .\next_auto_state_8__N_1686[7] (next_auto_state_8__N_1686[7]), 
            .n52359(n52359), .\swa_swb_val[1] (swa_swb_val[1])) /* synthesis syn_module_defined=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(281[17] 287[6])
    pwm_generator pwm_generator (.us_clk(us_clk), .us_clk_enable_61(us_clk_enable_61), 
            .high_counter_9__N_4408(high_counter_9__N_4408), .\next_state_2__N_4443[0] (next_state_2__N_4443[0]), 
            .GND_net(GND_net), .n53885(n53885), .resetn(resetn), .motor_4_pwm_c(motor_4_pwm_c), 
            .motor_3_pwm_c(motor_3_pwm_c), .motor_2_pwm_c(motor_2_pwm_c), 
            .motor_1_pwm_c(motor_1_pwm_c)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(495[19] 507[25])
    yaw_angle_accumulator YAAc (.n52179(n52179), .\state[5] (state_adj_5499[5]), 
            .\state[6] (state_adj_5499[6]), .n27995(n27995), .n37479(n37479)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(397[28] 413[10])
    \uart_top(NUM_DEBUG_ELEMENTS=8'b010010,FIXED_INTERVAL=0)  uart (.\tx_byte_index[0] (tx_byte_index[0]), 
            .\tx_byte_index[1] (tx_byte_index[1]), .n44797(n44797), .swa_swb_val({swa_swb_val}), 
            .n52359(n52359), .\led_data[0] (led_data[0]), .\led_data[3] (led_data[3]), 
            .\led_data[2] (led_data[2]), .\led_data[1] (led_data[1]), .n50(n50), 
            .n52(n52), .VL53L1X_chip_id({VL53L1X_chip_id}), .n43303(n43303), 
            .n43217(n43217), .\state[2] (state_adj_5499[2]), .n41683(n41683), 
            .\amc_debug[6] (amc_debug[6]), .\amc_debug[5] (amc_debug[5]), 
            .\state[5] (state_adj_5499[5]), .n52341(n52341), .n52342(n52342), 
            .latched_pitch({latched_pitch}), .n15182(n15182), .\z_linear_velocity[10] (z_linear_velocity[10]), 
            .\z_linear_velocity[8] (z_linear_velocity[8]), .\z_linear_velocity[9] (z_linear_velocity[9]), 
            .\z_linear_velocity[11] (z_linear_velocity[11]), .sys_clk(sys_clk), 
            .\next_state[0] (next_state_adj_5498[0]), .\tx_word_index[1] (tx_word_index[1]), 
            .VL53L1X_firm_rdy({VL53L1X_firm_rdy}), .throttle_val({throttle_val}), 
            .n49177(n49177), .\amc_debug[3] (amc_debug[3]), .\amc_debug[2] (amc_debug[2]), 
            .\amc_debug[1] (amc_debug[1]), .\amc_debug[7] (amc_debug[7]), 
            .\VL53L1X_range_mm[9] (VL53L1X_range_mm[9]), .\VL53L1X_range_mm[11] (VL53L1X_range_mm[11]), 
            .\VL53L1X_range_mm[10] (VL53L1X_range_mm[10]), .\VL53L1X_range_mm[15] (VL53L1X_range_mm[15]), 
            .\VL53L1X_range_mm[14] (VL53L1X_range_mm[14]), .\VL53L1X_range_mm[13] (VL53L1X_range_mm[13]), 
            .\z_linear_velocity[13] (z_linear_velocity[13]), .\z_linear_velocity[15] (z_linear_velocity[15]), 
            .\z_linear_velocity[14] (z_linear_velocity[14]), .n48813(n48813), 
            .n52441(n52441), .n52456(n52456), .yaw_val({yaw_val}), .n34690(n34690), 
            .n34692(n34692), .\latched_roll[2] (latched_roll[2]), .\state[6] (state_adj_5499[6]), 
            .\VL53L1X_range_mm[4] (VL53L1X_range_mm[4]), .\VL53L1X_range_mm[7] (VL53L1X_range_mm[7]), 
            .\VL53L1X_range_mm[6] (VL53L1X_range_mm[6]), .\VL53L1X_range_mm[5] (VL53L1X_range_mm[5]), 
            .n43332(n43332), .n43302(n43302), .\z_linear_velocity[7] (z_linear_velocity[7]), 
            .\z_linear_velocity[4] (z_linear_velocity[4]), .\z_linear_velocity[6] (z_linear_velocity[6]), 
            .\z_linear_velocity[5] (z_linear_velocity[5]), .\latched_roll[5] (latched_roll[5]), 
            .\latched_roll[7] (latched_roll[7]), .\latched_roll[6] (latched_roll[6]), 
            .\VL53L1X_range_mm[12] (VL53L1X_range_mm[12]), .\z_linear_velocity[12] (z_linear_velocity[12]), 
            .n44(n44), .n37479(n37479), .\led_data[4] (led_data[4]), .n52179(n52179), 
            .n37731(n37731), .n1406(n1406), .n27995(n27995), .n38(n38), 
            .\z_linear_velocity[3] (z_linear_velocity[3]), .\z_linear_velocity[2] (z_linear_velocity[2]), 
            .\z_linear_velocity[1] (z_linear_velocity[1]), .n34474(n34474), 
            .VL53L1X_data_rdy({VL53L1X_data_rdy}), .n43386(n43386), .n34665(n34665), 
            .n51335(n51335), .\latched_roll[4] (latched_roll[4]), .\amc_debug[4] (amc_debug[4]), 
            .\amc_debug[8] (amc_debug[8]), .n48820(n48820), .GND_net(GND_net), 
            .n52092(n52092), .n27(n27), .resetn_derived_2(resetn_derived_2), 
            .n51271(n51271), .n51272(n51272), .n43221(n43221), .n43225(n43225), 
            .n10(n10), .\amc_debug[0] (amc_debug[0]), .n43309(n43309), 
            .n48081(n48081), .n48828(n48828), .n49185(n49185), .n52267(n52267), 
            .n52328(n52328), .txrdy_n_c_7(txrdy_n_c_7), .n52255(n52255), 
            .n27734(n27734), .\VL53L1X_range_mm[8] (VL53L1X_range_mm[8]), 
            .n51044(n51044), .n52095(n52095), .n51041(n51041), .n123(n123), 
            .n43271(n43271), .n52390(n52390), .n51201(n51201), .n51202(n51202), 
            .n51159(n51159), .\i2c_device_driver_return_state[4] (i2c_device_driver_return_state[4]), 
            .n51273(n51273), .\VL53L1X_range_mm[1] (VL53L1X_range_mm[1]), 
            .\VL53L1X_range_mm[2] (VL53L1X_range_mm[2]), .n52388(n52388), 
            .n52389(n52389), .n41688(n41688), .n52429(n52429), .n36752(n36752), 
            .n50674(n50674), .n51135(n51135), .n50715(n50715), .n25(n25), 
            .n64(n64), .\led_data_out_7__N_1[2] (led_data_out_7__N_1[2]), 
            .n50881(n50881), .n52168(n52168), .n52169(n52169), .\i2c_device_driver_return_state[0] (i2c_device_driver_return_state[0]), 
            .\i2c_device_driver_return_state[3] (i2c_device_driver_return_state[3]), 
            .n52457(n52457), .\next_dat_i_15__N_4452[3] (next_dat_i_15__N_4452[3]), 
            .\next_state_4__N_1567[2] (next_state_4__N_1567[2]), .sout_c(sout_c), 
            .sin_c(sin_c), .n53885(n53885), .rxrdy_n_c(rxrdy_n_c), .n53884(n53884)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(528[64] 562[6])
    FD1S3AX VL53L1X_range_mm_i0 (.D(next_VL53L1X_range_mm[0]), .CK(sys_clk), 
            .Q(VL53L1X_range_mm[0]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(612[14] 649[12])
    defparam VL53L1X_range_mm_i0.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module throttle_controller
//

module throttle_controller (\state[0] , us_clk, resetn_derived_2, state, 
            throttle_controller_active, resetn, n49522, \state[2]_adj_6 , 
            \next_state_14__N_2466[1] , n48787, n4, n52214, n8, n30695, 
            n8773, n67, amc_complete_signal, n37558, n39759, n52213, 
            next_state_4__N_1666, n52566, n38) /* synthesis syn_module_defined=1 */ ;
    output \state[0] ;
    input us_clk;
    input resetn_derived_2;
    input [4:0]state;
    output throttle_controller_active;
    input resetn;
    input n49522;
    output \state[2]_adj_6 ;
    input \next_state_14__N_2466[1] ;
    output n48787;
    input n4;
    output n52214;
    output n8;
    input n30695;
    output [0:0]n8773;
    output n67;
    input amc_complete_signal;
    input n37558;
    output n39759;
    input n52213;
    output next_state_4__N_1666;
    output n52566;
    input n38;
    
    wire us_clk /* synthesis SET_AS_NETWORK=us_clk, is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(221[10:16])
    wire [6:0]state_c;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/throttle_controller.v(51[15:20])
    
    wire n52247, n51784, n51781, n51786;
    wire [6:0]next_state_6__N_1958;
    
    wire n52565, n52564;
    wire [6:0]next_state_6__N_1980;
    
    wire n21596, n39751, n52181, n51782, n51783, n39786, n52461, 
        n52211, n39753, n39755, n20, n26707, n39700, n52415, n49265, 
        n49345, n52411, n52472, n52473, n52471, n49563, n52304;
    
    LUT4 i1_2_lut_rep_311_3_lut_4_lut (.A(state_c[1]), .B(state_c[6]), .C(state_c[5]), 
         .D(state_c[3]), .Z(n52247)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/throttle_controller.v(79[14] 81[12])
    defparam i1_2_lut_rep_311_3_lut_4_lut.init = 16'hfffe;
    LUT4 n51785_bdd_2_lut_4_lut (.A(n51784), .B(n51781), .C(state_c[3]), 
         .D(state_c[6]), .Z(n51786)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam n51785_bdd_2_lut_4_lut.init = 16'hffca;
    FD1S3JX state_i0 (.D(next_state_6__N_1958[0]), .CK(us_clk), .PD(resetn_derived_2), 
            .Q(\state[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=25, LSE_LLINE=377, LSE_RLINE=389 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/throttle_controller.v(79[14] 81[12])
    defparam state_i0.GSR = "ENABLED";
    LUT4 n51048_bdd_2_lut_4_lut_then_4_lut (.A(state[0]), .B(state[1]), 
         .C(state[2]), .D(state[4]), .Z(n52565)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(74[31:36])
    defparam n51048_bdd_2_lut_4_lut_then_4_lut.init = 16'h0001;
    LUT4 n51048_bdd_2_lut_4_lut_else_4_lut (.A(state[0]), .B(state[1]), 
         .C(state[2]), .D(state[4]), .Z(n52564)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(74[31:36])
    defparam n51048_bdd_2_lut_4_lut_else_4_lut.init = 16'h0100;
    FD1P3AX active_signal_120 (.D(n49522), .SP(resetn), .CK(us_clk), .Q(throttle_controller_active)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=25, LSE_LLINE=377, LSE_RLINE=389 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/throttle_controller.v(136[14] 252[12])
    defparam active_signal_120.GSR = "DISABLED";
    FD1S3AX start_flag_110 (.D(n21596), .CK(us_clk), .Q(next_state_6__N_1980[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=25, LSE_LLINE=377, LSE_RLINE=389 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/throttle_controller.v(64[14] 71[42])
    defparam start_flag_110.GSR = "ENABLED";
    LUT4 i29135_4_lut_4_lut_4_lut (.A(state_c[1]), .B(state_c[6]), .C(state_c[3]), 
         .D(state_c[5]), .Z(n39751)) /* synthesis lut_function=(!(A+(B (C+(D))+!B (C (D)+!C !(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/throttle_controller.v(79[14] 81[12])
    defparam i29135_4_lut_4_lut_4_lut.init = 16'h0114;
    LUT4 i1_2_lut_rep_245_3_lut_4_lut (.A(\state[2]_adj_6 ), .B(n52247), 
         .C(\next_state_14__N_2466[1] ), .D(state_c[4]), .Z(n52181)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/throttle_controller.v(79[14] 81[12])
    defparam i1_2_lut_rep_245_3_lut_4_lut.init = 16'hfffe;
    LUT4 state_3__bdd_4_lut_40721 (.A(state_c[1]), .B(state_c[4]), .C(state_c[5]), 
         .D(\state[2]_adj_6 ), .Z(n51781)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam state_3__bdd_4_lut_40721.init = 16'hfffe;
    LUT4 state_1__bdd_4_lut_41233 (.A(state_c[4]), .B(state_c[5]), .C(next_state_6__N_1980[2]), 
         .D(\state[2]_adj_6 ), .Z(n51782)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;
    defparam state_1__bdd_4_lut_41233.init = 16'hffef;
    LUT4 state_1__bdd_3_lut (.A(state_c[4]), .B(state_c[5]), .C(\state[2]_adj_6 ), 
         .Z(n51783)) /* synthesis lut_function=(A (B+(C))+!A (B (C)+!B !(C))) */ ;
    defparam state_1__bdd_3_lut.init = 16'he9e9;
    LUT4 i29170_3_lut_4_lut_3_lut_4_lut (.A(state_c[1]), .B(state_c[6]), 
         .C(state_c[5]), .D(state_c[3]), .Z(n39786)) /* synthesis lut_function=(!(A+(B+(C (D)+!C !(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/throttle_controller.v(79[14] 81[12])
    defparam i29170_3_lut_4_lut_3_lut_4_lut.init = 16'h0110;
    LUT4 i111_3_lut_rep_278 (.A(n48787), .B(state[0]), .C(n4), .Z(n52214)) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(74[31:36])
    defparam i111_3_lut_rep_278.init = 16'ha8a8;
    LUT4 i19_4_lut_3_lut_4_lut (.A(state_c[3]), .B(n52461), .C(state_c[4]), 
         .D(state_c[5]), .Z(n8)) /* synthesis lut_function=(!(A+(B+(C (D)+!C !(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/throttle_controller.v(79[14] 81[12])
    defparam i19_4_lut_3_lut_4_lut.init = 16'h0110;
    LUT4 i1_2_lut_rep_275_3_lut_4_lut (.A(state_c[3]), .B(n52461), .C(\state[2]_adj_6 ), 
         .D(state_c[5]), .Z(n52211)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/throttle_controller.v(79[14] 81[12])
    defparam i1_2_lut_rep_275_3_lut_4_lut.init = 16'hfffe;
    LUT4 i29139_3_lut_4_lut (.A(state_c[4]), .B(n52211), .C(\state[0] ), 
         .D(n39753), .Z(n39755)) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/throttle_controller.v(79[14] 81[12])
    defparam i29139_3_lut_4_lut.init = 16'h1f10;
    FD1S3IX state_i5 (.D(n30695), .CK(us_clk), .CD(n20), .Q(state_c[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=25, LSE_LLINE=377, LSE_RLINE=389 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/throttle_controller.v(79[14] 81[12])
    defparam state_i5.GSR = "ENABLED";
    FD1S3IX state_i4 (.D(n26707), .CK(us_clk), .CD(\state[2]_adj_6 ), 
            .Q(state_c[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=25, LSE_LLINE=377, LSE_RLINE=389 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/throttle_controller.v(79[14] 81[12])
    defparam state_i4.GSR = "ENABLED";
    FD1S3IX state_i3 (.D(n26707), .CK(us_clk), .CD(n39700), .Q(state_c[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=25, LSE_LLINE=377, LSE_RLINE=389 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/throttle_controller.v(79[14] 81[12])
    defparam state_i3.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut (.A(state_c[4]), .B(n52211), .C(\state[0] ), 
         .D(\next_state_14__N_2466[1] ), .Z(next_state_6__N_1958[0])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/throttle_controller.v(79[14] 81[12])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0010;
    FD1S3IX state_i1 (.D(next_state_6__N_1958[1]), .CK(us_clk), .CD(resetn_derived_2), 
            .Q(state_c[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=25, LSE_LLINE=377, LSE_RLINE=389 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/throttle_controller.v(79[14] 81[12])
    defparam state_i1.GSR = "ENABLED";
    LUT4 i1_4_lut (.A(\state[0] ), .B(n39786), .C(n39753), .D(n52415), 
         .Z(n8773[0])) /* synthesis lut_function=(!(A+!(B (C+(D))+!B !((D)+!C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/throttle_controller.v(79[14] 81[12])
    defparam i1_4_lut.init = 16'h4450;
    LUT4 i5_4_lut (.A(n49265), .B(n49345), .C(state_c[1]), .D(n52411), 
         .Z(n67)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i5_4_lut.init = 16'h0010;
    LUT4 i38473_2_lut (.A(state_c[5]), .B(state_c[6]), .Z(n49265)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i38473_2_lut.init = 16'heeee;
    LUT4 i38550_2_lut (.A(\state[2]_adj_6 ), .B(state_c[3]), .Z(n49345)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i38550_2_lut.init = 16'heeee;
    LUT4 i1_3_lut (.A(n67), .B(amc_complete_signal), .C(next_state_6__N_1980[2]), 
         .Z(n21596)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/throttle_controller.v(51[15:20])
    defparam i1_3_lut.init = 16'hecec;
    LUT4 i29164_4_lut_4_lut_then_4_lut (.A(state_c[5]), .B(state_c[6]), 
         .C(state_c[1]), .D(\state[2]_adj_6 ), .Z(n52472)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/throttle_controller.v(79[14] 81[12])
    defparam i29164_4_lut_4_lut_then_4_lut.init = 16'h0001;
    LUT4 i106_2_lut_rep_475 (.A(\state[0] ), .B(state_c[4]), .Z(n52411)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i106_2_lut_rep_475.init = 16'heeee;
    LUT4 i2_3_lut_4_lut (.A(\state[0] ), .B(state_c[4]), .C(n52473), .D(resetn), 
         .Z(n26707)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;
    defparam i2_3_lut_4_lut.init = 16'h1000;
    PFUMX i40908 (.BLUT(n52471), .ALUT(n52472), .C0(state_c[3]), .Z(n52473));
    LUT4 i38746_2_lut_rep_479 (.A(state_c[4]), .B(\state[2]_adj_6 ), .Z(n52415)) /* synthesis lut_function=(!(A+(B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/throttle_controller.v(51[15:20])
    defparam i38746_2_lut_rep_479.init = 16'h1111;
    LUT4 i39798_2_lut_3_lut (.A(state_c[4]), .B(\state[2]_adj_6 ), .C(\state[0] ), 
         .Z(n49563)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/throttle_controller.v(51[15:20])
    defparam i39798_2_lut_3_lut.init = 16'hfefe;
    LUT4 i29164_4_lut_4_lut_else_4_lut (.A(state_c[5]), .B(state_c[6]), 
         .C(state_c[1]), .D(\state[2]_adj_6 ), .Z(n52471)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/throttle_controller.v(79[14] 81[12])
    defparam i29164_4_lut_4_lut_else_4_lut.init = 16'h0100;
    LUT4 i153_1_lut (.A(next_state_6__N_1980[2]), .Z(next_state_6__N_1980[1])) /* synthesis lut_function=(!(A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/throttle_controller.v(100[25:52])
    defparam i153_1_lut.init = 16'h5555;
    LUT4 i29158_1_lut (.A(state_c[4]), .Z(n20)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/throttle_controller.v(79[14] 81[12])
    defparam i29158_1_lut.init = 16'h5555;
    LUT4 i29084_1_lut (.A(\state[2]_adj_6 ), .Z(n39700)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/throttle_controller.v(79[14] 81[12])
    defparam i29084_1_lut.init = 16'h5555;
    LUT4 i29137_3_lut_3_lut_4_lut (.A(state_c[5]), .B(n52304), .C(state_c[4]), 
         .D(\state[2]_adj_6 ), .Z(n39753)) /* synthesis lut_function=(!(A+(B+(C (D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/throttle_controller.v(79[14] 81[12])
    defparam i29137_3_lut_3_lut_4_lut.init = 16'h0111;
    LUT4 i2_4_lut (.A(state[3]), .B(state[2]), .C(state[0]), .D(n37558), 
         .Z(n48787)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+((D)+!C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(74[31:36])
    defparam i2_4_lut.init = 16'hffed;
    PFUMX i40669 (.BLUT(n51786), .ALUT(n52181), .C0(\state[0] ), .Z(next_state_6__N_1958[1]));
    PFUMX i40667 (.BLUT(n51783), .ALUT(n51782), .C0(state_c[1]), .Z(n51784));
    PFUMX i29143 (.BLUT(n39751), .ALUT(n39755), .C0(n49563), .Z(n39759));
    LUT4 i3_4_lut (.A(state[0]), .B(n52214), .C(n52213), .D(\next_state_14__N_2466[1] ), 
         .Z(next_state_4__N_1666)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i3_4_lut.init = 16'h0020;
    PFUMX i40970 (.BLUT(n52564), .ALUT(n52565), .C0(state[3]), .Z(n52566));
    LUT4 i1_2_lut_rep_525 (.A(state_c[1]), .B(state_c[6]), .Z(n52461)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/throttle_controller.v(79[14] 81[12])
    defparam i1_2_lut_rep_525.init = 16'heeee;
    FD1S3IX state_i2 (.D(n38), .CK(us_clk), .CD(next_state_6__N_1980[1]), 
            .Q(\state[2]_adj_6 )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=25, LSE_LLINE=377, LSE_RLINE=389 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/throttle_controller.v(79[14] 81[12])
    defparam state_i2.GSR = "ENABLED";
    FD1S3IX state_i6 (.D(n30695), .CK(us_clk), .CD(state_c[4]), .Q(state_c[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=25, LSE_LLINE=377, LSE_RLINE=389 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/throttle_controller.v(79[14] 81[12])
    defparam state_i6.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_368_3_lut (.A(state_c[1]), .B(state_c[6]), .C(state_c[3]), 
         .Z(n52304)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/throttle_controller.v(79[14] 81[12])
    defparam i1_2_lut_rep_368_3_lut.init = 16'hfefe;
    
endmodule
//
// Verilog Description of module TSALL
// module not written out since it is a black-box. 
//

//
// Verilog Description of module PUR
// module not written out since it is a black-box. 
//

//
// Verilog Description of module us_clk
//

module us_clk (GND_net, us_clk, sys_clk) /* synthesis syn_module_defined=1 */ ;
    input GND_net;
    output us_clk;
    input sys_clk;
    
    wire us_clk /* synthesis SET_AS_NETWORK=us_clk, is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(221[10:16])
    wire sys_clk /* synthesis SET_AS_NETWORK=sys_clk, is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(220[10:17])
    
    wire n43776;
    wire [14:0]sys_clk_counter;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/us_clk.v(23[16:31])
    wire [14:0]n7;
    
    wire n43777, n16227, n43779, n43780, n30629;
    wire [14:0]sys_clk_counter_14__N_11;
    
    wire n43775, n29, n29_adj_5365, n27431, n6, n6_adj_5366, n15_adj_5367, 
        n20_adj_5368, n18_adj_5369, n43778, n43781;
    
    CCU2D add_7_5 (.A0(sys_clk_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(sys_clk_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43776), .COUT(n43777), .S0(n7[3]), .S1(n7[4]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/us_clk.v(39[32:54])
    defparam add_7_5.INIT0 = 16'h5aaa;
    defparam add_7_5.INIT1 = 16'h5aaa;
    defparam add_7_5.INJECT1_0 = "NO";
    defparam add_7_5.INJECT1_1 = "NO";
    FD1S3AY us_clk_16 (.D(n16227), .CK(sys_clk), .Q(us_clk)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=25, LSE_LLINE=249, LSE_RLINE=252 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/us_clk.v(30[14] 39[55])
    defparam us_clk_16.GSR = "ENABLED";
    CCU2D add_7_11 (.A0(sys_clk_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(sys_clk_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43779), .COUT(n43780), .S0(n7[9]), .S1(n7[10]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/us_clk.v(39[32:54])
    defparam add_7_11.INIT0 = 16'h5aaa;
    defparam add_7_11.INIT1 = 16'h5aaa;
    defparam add_7_11.INJECT1_0 = "NO";
    defparam add_7_11.INJECT1_1 = "NO";
    FD1S3IX sys_clk_counter_i14 (.D(n7[14]), .CK(sys_clk), .CD(n30629), 
            .Q(sys_clk_counter[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=25, LSE_LLINE=249, LSE_RLINE=252 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/us_clk.v(30[14] 39[55])
    defparam sys_clk_counter_i14.GSR = "ENABLED";
    FD1S3IX sys_clk_counter_i13 (.D(n7[13]), .CK(sys_clk), .CD(n30629), 
            .Q(sys_clk_counter[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=25, LSE_LLINE=249, LSE_RLINE=252 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/us_clk.v(30[14] 39[55])
    defparam sys_clk_counter_i13.GSR = "ENABLED";
    FD1S3IX sys_clk_counter_i12 (.D(n7[12]), .CK(sys_clk), .CD(n30629), 
            .Q(sys_clk_counter[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=25, LSE_LLINE=249, LSE_RLINE=252 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/us_clk.v(30[14] 39[55])
    defparam sys_clk_counter_i12.GSR = "ENABLED";
    FD1S3IX sys_clk_counter_i11 (.D(n7[11]), .CK(sys_clk), .CD(n30629), 
            .Q(sys_clk_counter[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=25, LSE_LLINE=249, LSE_RLINE=252 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/us_clk.v(30[14] 39[55])
    defparam sys_clk_counter_i11.GSR = "ENABLED";
    FD1S3IX sys_clk_counter_i10 (.D(n7[10]), .CK(sys_clk), .CD(n30629), 
            .Q(sys_clk_counter[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=25, LSE_LLINE=249, LSE_RLINE=252 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/us_clk.v(30[14] 39[55])
    defparam sys_clk_counter_i10.GSR = "ENABLED";
    FD1S3IX sys_clk_counter_i9 (.D(n7[9]), .CK(sys_clk), .CD(n30629), 
            .Q(sys_clk_counter[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=25, LSE_LLINE=249, LSE_RLINE=252 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/us_clk.v(30[14] 39[55])
    defparam sys_clk_counter_i9.GSR = "ENABLED";
    FD1S3IX sys_clk_counter_i8 (.D(n7[8]), .CK(sys_clk), .CD(n30629), 
            .Q(sys_clk_counter[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=25, LSE_LLINE=249, LSE_RLINE=252 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/us_clk.v(30[14] 39[55])
    defparam sys_clk_counter_i8.GSR = "ENABLED";
    FD1S3IX sys_clk_counter_i7 (.D(n7[7]), .CK(sys_clk), .CD(n30629), 
            .Q(sys_clk_counter[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=25, LSE_LLINE=249, LSE_RLINE=252 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/us_clk.v(30[14] 39[55])
    defparam sys_clk_counter_i7.GSR = "ENABLED";
    FD1S3IX sys_clk_counter_i6 (.D(n7[6]), .CK(sys_clk), .CD(n30629), 
            .Q(sys_clk_counter[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=25, LSE_LLINE=249, LSE_RLINE=252 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/us_clk.v(30[14] 39[55])
    defparam sys_clk_counter_i6.GSR = "ENABLED";
    FD1S3IX sys_clk_counter_i5 (.D(n7[5]), .CK(sys_clk), .CD(n30629), 
            .Q(sys_clk_counter[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=25, LSE_LLINE=249, LSE_RLINE=252 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/us_clk.v(30[14] 39[55])
    defparam sys_clk_counter_i5.GSR = "ENABLED";
    FD1S3IX sys_clk_counter_i3 (.D(n7[3]), .CK(sys_clk), .CD(n30629), 
            .Q(sys_clk_counter[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=25, LSE_LLINE=249, LSE_RLINE=252 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/us_clk.v(30[14] 39[55])
    defparam sys_clk_counter_i3.GSR = "ENABLED";
    FD1S3AX sys_clk_counter_i2 (.D(sys_clk_counter_14__N_11[2]), .CK(sys_clk), 
            .Q(sys_clk_counter[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=25, LSE_LLINE=249, LSE_RLINE=252 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/us_clk.v(30[14] 39[55])
    defparam sys_clk_counter_i2.GSR = "ENABLED";
    FD1S3IX sys_clk_counter_i1 (.D(n7[1]), .CK(sys_clk), .CD(n30629), 
            .Q(sys_clk_counter[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=25, LSE_LLINE=249, LSE_RLINE=252 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/us_clk.v(30[14] 39[55])
    defparam sys_clk_counter_i1.GSR = "ENABLED";
    CCU2D add_7_3 (.A0(sys_clk_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(sys_clk_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43775), .COUT(n43776), .S0(n7[1]), .S1(n7[2]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/us_clk.v(39[32:54])
    defparam add_7_3.INIT0 = 16'h5aaa;
    defparam add_7_3.INIT1 = 16'h5aaa;
    defparam add_7_3.INJECT1_0 = "NO";
    defparam add_7_3.INJECT1_1 = "NO";
    LUT4 i25759_3_lut (.A(us_clk), .B(n29), .C(n29_adj_5365), .Z(n16227)) /* synthesis lut_function=(A (B)+!A !((C)+!B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/us_clk.v(30[14] 39[55])
    defparam i25759_3_lut.init = 16'h8c8c;
    LUT4 i4_4_lut (.A(sys_clk_counter[1]), .B(sys_clk_counter[4]), .C(n27431), 
         .D(n6), .Z(n29)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i4_4_lut.init = 16'hfff7;
    LUT4 i1_2_lut (.A(sys_clk_counter[5]), .B(sys_clk_counter[2]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i4_4_lut_adj_515 (.A(sys_clk_counter[2]), .B(sys_clk_counter[5]), 
         .C(n27431), .D(n6_adj_5366), .Z(n29_adj_5365)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;
    defparam i4_4_lut_adj_515.init = 16'hfff7;
    LUT4 i1_2_lut_adj_516 (.A(sys_clk_counter[4]), .B(sys_clk_counter[1]), 
         .Z(n6_adj_5366)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_516.init = 16'heeee;
    LUT4 i10_4_lut (.A(n15_adj_5367), .B(n20_adj_5368), .C(sys_clk_counter[0]), 
         .D(sys_clk_counter[12]), .Z(n27431)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/us_clk.v(34[18:55])
    defparam i10_4_lut.init = 16'hffef;
    LUT4 i4_2_lut (.A(sys_clk_counter[7]), .B(sys_clk_counter[9]), .Z(n15_adj_5367)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/us_clk.v(34[18:55])
    defparam i4_2_lut.init = 16'heeee;
    LUT4 i9_4_lut (.A(sys_clk_counter[14]), .B(n18_adj_5369), .C(sys_clk_counter[6]), 
         .D(sys_clk_counter[8]), .Z(n20_adj_5368)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/us_clk.v(34[18:55])
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 i7_4_lut (.A(sys_clk_counter[10]), .B(sys_clk_counter[3]), .C(sys_clk_counter[11]), 
         .D(sys_clk_counter[13]), .Z(n18_adj_5369)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/us_clk.v(34[18:55])
    defparam i7_4_lut.init = 16'hfffe;
    LUT4 i26393_3_lut (.A(n7[4]), .B(n29), .C(n29_adj_5365), .Z(sys_clk_counter_14__N_11[4])) /* synthesis lut_function=(A ((C)+!B)+!A !(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/us_clk.v(34[14] 39[55])
    defparam i26393_3_lut.init = 16'hb3b3;
    CCU2D add_7_9 (.A0(sys_clk_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(sys_clk_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43778), .COUT(n43779), .S0(n7[7]), .S1(n7[8]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/us_clk.v(39[32:54])
    defparam add_7_9.INIT0 = 16'h5aaa;
    defparam add_7_9.INIT1 = 16'h5aaa;
    defparam add_7_9.INJECT1_0 = "NO";
    defparam add_7_9.INJECT1_1 = "NO";
    CCU2D add_7_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(sys_clk_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n43775), .S1(n7[0]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/us_clk.v(39[32:54])
    defparam add_7_1.INIT0 = 16'hF000;
    defparam add_7_1.INIT1 = 16'h5555;
    defparam add_7_1.INJECT1_0 = "NO";
    defparam add_7_1.INJECT1_1 = "NO";
    CCU2D add_7_15 (.A0(sys_clk_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(sys_clk_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43781), .S0(n7[13]), .S1(n7[14]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/us_clk.v(39[32:54])
    defparam add_7_15.INIT0 = 16'h5aaa;
    defparam add_7_15.INIT1 = 16'h5aaa;
    defparam add_7_15.INJECT1_0 = "NO";
    defparam add_7_15.INJECT1_1 = "NO";
    CCU2D add_7_13 (.A0(sys_clk_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(sys_clk_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43780), .COUT(n43781), .S0(n7[11]), .S1(n7[12]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/us_clk.v(39[32:54])
    defparam add_7_13.INIT0 = 16'h5aaa;
    defparam add_7_13.INIT1 = 16'h5aaa;
    defparam add_7_13.INJECT1_0 = "NO";
    defparam add_7_13.INJECT1_1 = "NO";
    LUT4 i39434_2_lut (.A(n29_adj_5365), .B(n29), .Z(n30629)) /* synthesis lut_function=(!(A (B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/us_clk.v(34[14] 39[55])
    defparam i39434_2_lut.init = 16'h7777;
    LUT4 i26400_3_lut (.A(n7[2]), .B(n29), .C(n29_adj_5365), .Z(sys_clk_counter_14__N_11[2])) /* synthesis lut_function=(A ((C)+!B)+!A !(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/us_clk.v(34[14] 39[55])
    defparam i26400_3_lut.init = 16'hb3b3;
    CCU2D add_7_7 (.A0(sys_clk_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(sys_clk_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43777), .COUT(n43778), .S0(n7[5]), .S1(n7[6]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/us_clk.v(39[32:54])
    defparam add_7_7.INIT0 = 16'h5aaa;
    defparam add_7_7.INIT1 = 16'h5aaa;
    defparam add_7_7.INJECT1_0 = "NO";
    defparam add_7_7.INJECT1_1 = "NO";
    FD1S3AX sys_clk_counter_i4 (.D(sys_clk_counter_14__N_11[4]), .CK(sys_clk), 
            .Q(sys_clk_counter[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=25, LSE_LLINE=249, LSE_RLINE=252 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/us_clk.v(30[14] 39[55])
    defparam sys_clk_counter_i4.GSR = "ENABLED";
    FD1S3IX sys_clk_counter_i0 (.D(n7[0]), .CK(sys_clk), .CD(n30629), 
            .Q(sys_clk_counter[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=12, LSE_RCOL=25, LSE_LLINE=249, LSE_RLINE=252 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/us_clk.v(30[14] 39[55])
    defparam sys_clk_counter_i0.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module receiver
//

module receiver (state_2__N_199_c_1, us_clk, GND_net, yaw_val, n43271, 
            n52456, n51041, state_2__N_84_c_1, resetn, resetn_derived_2, 
            \i2c_top_debug[1] , n52306, wd_event_active, n52205, n44, 
            n44797, n64, \next_state[0] , n33315, count__auto_time_ms_27__N_1639, 
            n52318, n52142, \i2c_top_debug[5] , byte_rd_left_5__N_1255, 
            throttle_val, n52441, n51044, n52429, swa_swb_val, state_2__N_199_c_1_adj_2, 
            state_2__N_199_c_1_adj_3, \latched_roll[7] , \latched_roll[6] , 
            \latched_roll[5] , \latched_roll[4] , \latched_roll[2] , n48820, 
            state_2__N_199_c_1_adj_4, n1406, latched_pitch, n52328, 
            \tx_byte_index[0] , n52095, n27, \tx_byte_index[1] , \tx_word_index[1] , 
            n36649, n34665, n51272, n51271, n51273, n51202, n51159, 
            n51201, n34692, n36752, n34690) /* synthesis syn_module_defined=1 */ ;
    input state_2__N_199_c_1;
    input us_clk;
    input GND_net;
    output [7:0]yaw_val;
    output n43271;
    output n52456;
    output n51041;
    input state_2__N_84_c_1;
    input resetn;
    output resetn_derived_2;
    input \i2c_top_debug[1] ;
    input n52306;
    input wd_event_active;
    output n52205;
    input n44;
    input n44797;
    input n64;
    output \next_state[0] ;
    input n33315;
    output count__auto_time_ms_27__N_1639;
    output n52318;
    input n52142;
    input \i2c_top_debug[5] ;
    output byte_rd_left_5__N_1255;
    output [7:0]throttle_val;
    output n52441;
    output n51044;
    output n52429;
    output [7:0]swa_swb_val;
    input state_2__N_199_c_1_adj_2;
    input state_2__N_199_c_1_adj_3;
    output \latched_roll[7] ;
    output \latched_roll[6] ;
    output \latched_roll[5] ;
    output \latched_roll[4] ;
    output \latched_roll[2] ;
    output n48820;
    input state_2__N_199_c_1_adj_4;
    output n1406;
    output [7:0]latched_pitch;
    input n52328;
    input \tx_byte_index[0] ;
    output n52095;
    output n27;
    input \tx_byte_index[1] ;
    input \tx_word_index[1] ;
    input n36649;
    output n34665;
    input n51272;
    input n51271;
    output n51273;
    output n51202;
    output n51159;
    output n51201;
    output n34692;
    output n36752;
    output n34690;
    
    wire us_clk /* synthesis SET_AS_NETWORK=us_clk, is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(221[10:16])
    wire [15:0]yaw_pwm_pulse_length_us;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/receiver.v(52[9:32])
    wire [15:0]throttle_pwm_pulse_length_us;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/receiver.v(51[9:37])
    wire [15:0]swa_swb_pwm_pulse_length_us;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/receiver.v(57[9:36])
    wire [15:0]roll_pwm_pulse_length_us;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/receiver.v(53[9:33])
    wire [7:0]latched_roll;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/angle_controller.v(84[74:86])
    wire [15:0]pitch_pwm_pulse_length_us;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/receiver.v(54[9:34])
    
    pwm_reader yaw_reader (.state_2__N_199_c_1(state_2__N_199_c_1), .us_clk(us_clk), 
            .GND_net(GND_net), .\yaw_pwm_pulse_length_us[2] (yaw_pwm_pulse_length_us[2]), 
            .\yaw_pwm_pulse_length_us[3] (yaw_pwm_pulse_length_us[3]), .\yaw_pwm_pulse_length_us[4] (yaw_pwm_pulse_length_us[4]), 
            .\yaw_pwm_pulse_length_us[5] (yaw_pwm_pulse_length_us[5]), .\yaw_pwm_pulse_length_us[6] (yaw_pwm_pulse_length_us[6]), 
            .\yaw_pwm_pulse_length_us[7] (yaw_pwm_pulse_length_us[7]), .\yaw_pwm_pulse_length_us[8] (yaw_pwm_pulse_length_us[8]), 
            .\yaw_pwm_pulse_length_us[9] (yaw_pwm_pulse_length_us[9])) /* synthesis syn_module_defined=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/receiver.v(76[51] 82[25])
    pwm_to_value yaw_pwm_to_value (.yaw_val({yaw_val}), .us_clk(us_clk), 
            .\yaw_pwm_pulse_length_us[2] (yaw_pwm_pulse_length_us[2]), .\yaw_pwm_pulse_length_us[5] (yaw_pwm_pulse_length_us[5]), 
            .\yaw_pwm_pulse_length_us[7] (yaw_pwm_pulse_length_us[7]), .\yaw_pwm_pulse_length_us[6] (yaw_pwm_pulse_length_us[6]), 
            .\yaw_pwm_pulse_length_us[8] (yaw_pwm_pulse_length_us[8]), .\yaw_pwm_pulse_length_us[4] (yaw_pwm_pulse_length_us[4]), 
            .\yaw_pwm_pulse_length_us[3] (yaw_pwm_pulse_length_us[3]), .\yaw_pwm_pulse_length_us[9] (yaw_pwm_pulse_length_us[9]), 
            .n43271(n43271), .n52456(n52456), .n51041(n51041)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/receiver.v(84[18] 89[25])
    \pwm_reader(DEFAULT_PWM_TIME_HIGH_US=16'b01111101000)  throttle_reader (.state_2__N_84_c_1(state_2__N_84_c_1), 
            .GND_net(GND_net), .us_clk(us_clk), .resetn(resetn), .resetn_derived_2(resetn_derived_2), 
            .\i2c_top_debug[1] (\i2c_top_debug[1] ), .n52306(n52306), .wd_event_active(wd_event_active), 
            .n52205(n52205), .n44(n44), .n44797(n44797), .n64(n64), 
            .\next_state[0] (\next_state[0] ), .n33315(n33315), .count__auto_time_ms_27__N_1639(count__auto_time_ms_27__N_1639), 
            .n52318(n52318), .n52142(n52142), .\i2c_top_debug[5] (\i2c_top_debug[5] ), 
            .byte_rd_left_5__N_1255(byte_rd_left_5__N_1255), .\throttle_pwm_pulse_length_us[4] (throttle_pwm_pulse_length_us[4]), 
            .\throttle_pwm_pulse_length_us[9] (throttle_pwm_pulse_length_us[9]), 
            .\throttle_pwm_pulse_length_us[8] (throttle_pwm_pulse_length_us[8]), 
            .\throttle_pwm_pulse_length_us[7] (throttle_pwm_pulse_length_us[7]), 
            .\throttle_pwm_pulse_length_us[6] (throttle_pwm_pulse_length_us[6]), 
            .\throttle_pwm_pulse_length_us[5] (throttle_pwm_pulse_length_us[5]), 
            .\throttle_pwm_pulse_length_us[3] (throttle_pwm_pulse_length_us[3]), 
            .\throttle_pwm_pulse_length_us[2] (throttle_pwm_pulse_length_us[2])) /* synthesis syn_module_defined=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/receiver.v(60[56] 66[25])
    pwm_to_value_U0 throttle_pwm_to_value (.throttle_val({throttle_val}), 
            .us_clk(us_clk), .\throttle_pwm_pulse_length_us[2] (throttle_pwm_pulse_length_us[2]), 
            .\throttle_pwm_pulse_length_us[5] (throttle_pwm_pulse_length_us[5]), 
            .\throttle_pwm_pulse_length_us[7] (throttle_pwm_pulse_length_us[7]), 
            .\throttle_pwm_pulse_length_us[6] (throttle_pwm_pulse_length_us[6]), 
            .\throttle_pwm_pulse_length_us[8] (throttle_pwm_pulse_length_us[8]), 
            .n52441(n52441), .n51044(n51044), .\throttle_pwm_pulse_length_us[9] (throttle_pwm_pulse_length_us[9]), 
            .\throttle_pwm_pulse_length_us[4] (throttle_pwm_pulse_length_us[4]), 
            .\throttle_pwm_pulse_length_us[3] (throttle_pwm_pulse_length_us[3]), 
            .n52429(n52429)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/receiver.v(68[18] 73[25])
    pwm_to_value_U1 swab_pwm_to_value (.\swa_swb_pwm_pulse_length_us[5] (swa_swb_pwm_pulse_length_us[5]), 
            .\swa_swb_pwm_pulse_length_us[7] (swa_swb_pwm_pulse_length_us[7]), 
            .\swa_swb_pwm_pulse_length_us[6] (swa_swb_pwm_pulse_length_us[6]), 
            .swa_swb_val({swa_swb_val}), .us_clk(us_clk), .\swa_swb_pwm_pulse_length_us[2] (swa_swb_pwm_pulse_length_us[2]), 
            .\swa_swb_pwm_pulse_length_us[8] (swa_swb_pwm_pulse_length_us[8]), 
            .\swa_swb_pwm_pulse_length_us[9] (swa_swb_pwm_pulse_length_us[9]), 
            .\swa_swb_pwm_pulse_length_us[4] (swa_swb_pwm_pulse_length_us[4]), 
            .\swa_swb_pwm_pulse_length_us[3] (swa_swb_pwm_pulse_length_us[3])) /* synthesis syn_module_defined=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/receiver.v(167[18] 172[25])
    pwm_reader_U2 swa_swb_reader (.state_2__N_199_c_1(state_2__N_199_c_1_adj_2), 
            .us_clk(us_clk), .GND_net(GND_net), .\swa_swb_pwm_pulse_length_us[2] (swa_swb_pwm_pulse_length_us[2]), 
            .\swa_swb_pwm_pulse_length_us[3] (swa_swb_pwm_pulse_length_us[3]), 
            .\swa_swb_pwm_pulse_length_us[4] (swa_swb_pwm_pulse_length_us[4]), 
            .\swa_swb_pwm_pulse_length_us[5] (swa_swb_pwm_pulse_length_us[5]), 
            .\swa_swb_pwm_pulse_length_us[6] (swa_swb_pwm_pulse_length_us[6]), 
            .\swa_swb_pwm_pulse_length_us[7] (swa_swb_pwm_pulse_length_us[7]), 
            .\swa_swb_pwm_pulse_length_us[8] (swa_swb_pwm_pulse_length_us[8]), 
            .\swa_swb_pwm_pulse_length_us[9] (swa_swb_pwm_pulse_length_us[9])) /* synthesis syn_module_defined=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/receiver.v(159[5] 165[25])
    pwm_reader_U3 roll_reader (.state_2__N_199_c_1(state_2__N_199_c_1_adj_3), 
            .us_clk(us_clk), .GND_net(GND_net), .\roll_pwm_pulse_length_us[2] (roll_pwm_pulse_length_us[2]), 
            .\roll_pwm_pulse_length_us[3] (roll_pwm_pulse_length_us[3]), .\roll_pwm_pulse_length_us[4] (roll_pwm_pulse_length_us[4]), 
            .\roll_pwm_pulse_length_us[5] (roll_pwm_pulse_length_us[5]), .\roll_pwm_pulse_length_us[6] (roll_pwm_pulse_length_us[6]), 
            .\roll_pwm_pulse_length_us[7] (roll_pwm_pulse_length_us[7]), .\roll_pwm_pulse_length_us[8] (roll_pwm_pulse_length_us[8]), 
            .\roll_pwm_pulse_length_us[9] (roll_pwm_pulse_length_us[9])) /* synthesis syn_module_defined=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/receiver.v(92[52] 98[25])
    pwm_to_value_U4 roll_pwm_to_value (.latched_roll({\latched_roll[7] , \latched_roll[6] , 
            \latched_roll[5] , \latched_roll[4] , latched_roll[3], \latched_roll[2] , 
            latched_roll[1:0]}), .us_clk(us_clk), .\roll_pwm_pulse_length_us[2] (roll_pwm_pulse_length_us[2]), 
            .\roll_pwm_pulse_length_us[5] (roll_pwm_pulse_length_us[5]), .\roll_pwm_pulse_length_us[7] (roll_pwm_pulse_length_us[7]), 
            .\roll_pwm_pulse_length_us[6] (roll_pwm_pulse_length_us[6]), .\roll_pwm_pulse_length_us[4] (roll_pwm_pulse_length_us[4]), 
            .\roll_pwm_pulse_length_us[3] (roll_pwm_pulse_length_us[3]), .\roll_pwm_pulse_length_us[8] (roll_pwm_pulse_length_us[8]), 
            .n48820(n48820), .\roll_pwm_pulse_length_us[9] (roll_pwm_pulse_length_us[9])) /* synthesis syn_module_defined=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/receiver.v(100[18] 105[25])
    pwm_reader_U5 pitch_reader (.state_2__N_199_c_1(state_2__N_199_c_1_adj_4), 
            .us_clk(us_clk), .GND_net(GND_net), .\pitch_pwm_pulse_length_us[2] (pitch_pwm_pulse_length_us[2]), 
            .\pitch_pwm_pulse_length_us[3] (pitch_pwm_pulse_length_us[3]), 
            .\pitch_pwm_pulse_length_us[4] (pitch_pwm_pulse_length_us[4]), 
            .\pitch_pwm_pulse_length_us[5] (pitch_pwm_pulse_length_us[5]), 
            .\pitch_pwm_pulse_length_us[6] (pitch_pwm_pulse_length_us[6]), 
            .\pitch_pwm_pulse_length_us[7] (pitch_pwm_pulse_length_us[7]), 
            .\pitch_pwm_pulse_length_us[8] (pitch_pwm_pulse_length_us[8]), 
            .\pitch_pwm_pulse_length_us[9] (pitch_pwm_pulse_length_us[9])) /* synthesis syn_module_defined=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/receiver.v(108[53] 114[25])
    pwm_to_value_U6 pitch_pwm_to_value (.\latched_roll[2] (\latched_roll[2] ), 
            .\latched_roll[3] (latched_roll[3]), .\latched_roll[1] (latched_roll[1]), 
            .n1406(n1406), .latched_pitch({latched_pitch}), .us_clk(us_clk), 
            .\pitch_pwm_pulse_length_us[2] (pitch_pwm_pulse_length_us[2]), 
            .n52328(n52328), .\tx_byte_index[0] (\tx_byte_index[0] ), .n52095(n52095), 
            .n27(n27), .\tx_byte_index[1] (\tx_byte_index[1] ), .\tx_word_index[1] (\tx_word_index[1] ), 
            .n36649(n36649), .n34665(n34665), .\pitch_pwm_pulse_length_us[5] (pitch_pwm_pulse_length_us[5]), 
            .\pitch_pwm_pulse_length_us[7] (pitch_pwm_pulse_length_us[7]), 
            .\pitch_pwm_pulse_length_us[6] (pitch_pwm_pulse_length_us[6]), 
            .\pitch_pwm_pulse_length_us[4] (pitch_pwm_pulse_length_us[4]), 
            .\pitch_pwm_pulse_length_us[3] (pitch_pwm_pulse_length_us[3]), 
            .n51272(n51272), .n51271(n51271), .n51273(n51273), .\latched_roll[0] (latched_roll[0]), 
            .n51202(n51202), .n51159(n51159), .\swa_swb_val[0] (swa_swb_val[0]), 
            .\swa_swb_val[1] (swa_swb_val[1]), .\swa_swb_val[2] (swa_swb_val[2]), 
            .\swa_swb_val[3] (swa_swb_val[3]), .n51201(n51201), .n34692(n34692), 
            .n36752(n36752), .\pitch_pwm_pulse_length_us[8] (pitch_pwm_pulse_length_us[8]), 
            .n34690(n34690), .\pitch_pwm_pulse_length_us[9] (pitch_pwm_pulse_length_us[9])) /* synthesis syn_module_defined=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/receiver.v(116[18] 121[25])
    
endmodule
//
// Verilog Description of module pwm_reader
//

module pwm_reader (state_2__N_199_c_1, us_clk, GND_net, \yaw_pwm_pulse_length_us[2] , 
            \yaw_pwm_pulse_length_us[3] , \yaw_pwm_pulse_length_us[4] , 
            \yaw_pwm_pulse_length_us[5] , \yaw_pwm_pulse_length_us[6] , 
            \yaw_pwm_pulse_length_us[7] , \yaw_pwm_pulse_length_us[8] , 
            \yaw_pwm_pulse_length_us[9] ) /* synthesis syn_module_defined=1 */ ;
    input state_2__N_199_c_1;
    input us_clk;
    input GND_net;
    output \yaw_pwm_pulse_length_us[2] ;
    output \yaw_pwm_pulse_length_us[3] ;
    output \yaw_pwm_pulse_length_us[4] ;
    output \yaw_pwm_pulse_length_us[5] ;
    output \yaw_pwm_pulse_length_us[6] ;
    output \yaw_pwm_pulse_length_us[7] ;
    output \yaw_pwm_pulse_length_us[8] ;
    output \yaw_pwm_pulse_length_us[9] ;
    
    wire us_clk /* synthesis SET_AS_NETWORK=us_clk, is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(221[10:16])
    wire [2:0]state;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(54[15:20])
    
    wire us_clk_enable_147;
    wire [15:0]time_high_count_15__N_224;
    wire [15:0]time_high_count_15__N_183;
    wire [15:0]time_high_count;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(57[16:31])
    
    wire us_clk_enable_56;
    wire [2:0]state_2__N_180;
    
    wire n52458, n62, n80, n152, n35595, n8, n4, n35593, n4_adj_5357, 
        pwm_pulse_level_flag, n46791, us_clk_enable_58, n50712, n50713, 
        n51068, n51067, n52394, n47221, n35569, n3, n51111, n51113, 
        n51110, n3_adj_5358, n51109, n3_adj_5359;
    wire [15:0]pwm_pulse_length_us_15__N_208;
    
    wire n7, n49525, n50714, n48052, n35596, n3_adj_5360, n3_adj_5361, 
        us_clk_enable_126, n36397, n46559, n43941, n43940, n43939, 
        n43938, n43937, n43936, n43935, n43934, n30688, n51115;
    
    LUT4 i20_4_lut_3_lut_4_lut (.A(state[1]), .B(state_2__N_199_c_1), .C(state[0]), 
         .D(state[2]), .Z(us_clk_enable_147)) /* synthesis lut_function=(A (B ((D)+!C)+!B (D))+!A !(D)) */ ;
    defparam i20_4_lut_3_lut_4_lut.init = 16'haa5d;
    LUT4 i1_2_lut_4_lut (.A(state[2]), .B(state[1]), .C(state[0]), .D(time_high_count_15__N_224[1]), 
         .Z(time_high_count_15__N_183[1])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h0400;
    FD1P3AX time_high_count_i0 (.D(time_high_count_15__N_183[0]), .SP(us_clk_enable_56), 
            .CK(us_clk), .Q(time_high_count[0])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=51, LSE_RCOL=25, LSE_LLINE=76, LSE_RLINE=82 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i0.GSR = "ENABLED";
    FD1S3AX state_i0 (.D(state_2__N_180[0]), .CK(us_clk), .Q(state[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=14, LSE_LCOL=51, LSE_RCOL=25, LSE_LLINE=76, LSE_RLINE=82 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam state_i0.GSR = "ENABLED";
    LUT4 i2_3_lut (.A(time_high_count[6]), .B(n52458), .C(time_high_count[10]), 
         .Z(n62)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(57[16:31])
    defparam i2_3_lut.init = 16'h8080;
    LUT4 i12_4_lut (.A(n80), .B(time_high_count[4]), .C(time_high_count[5]), 
         .D(n152), .Z(n35595)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A !(D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(57[16:31])
    defparam i12_4_lut.init = 16'h5700;
    LUT4 i24963_4_lut (.A(n152), .B(n8), .C(time_high_count[6]), .D(n4), 
         .Z(n35593)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(57[16:31])
    defparam i24963_4_lut.init = 16'hca0a;
    LUT4 i2_4_lut (.A(state[0]), .B(state_2__N_199_c_1), .C(state[1]), 
         .D(n4_adj_5357), .Z(us_clk_enable_56)) /* synthesis lut_function=((B (C)+!B (C+!(D)))+!A) */ ;
    defparam i2_4_lut.init = 16'hf5f7;
    LUT4 i1_2_lut (.A(state[2]), .B(pwm_pulse_level_flag), .Z(n4_adj_5357)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 state_2__N_199_c_1_bdd_4_lut_40214 (.A(state_2__N_199_c_1), .B(state[2]), 
         .C(state[0]), .D(state[1]), .Z(state_2__N_180[0])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B ((D)+!C)))) */ ;
    defparam state_2__N_199_c_1_bdd_4_lut_40214.init = 16'h3173;
    FD1S3IX state_i2 (.D(n46791), .CK(us_clk), .CD(state[2]), .Q(state[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=14, LSE_LCOL=51, LSE_RCOL=25, LSE_LLINE=76, LSE_RLINE=82 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam state_i2.GSR = "ENABLED";
    FD1S3AX state_i1 (.D(state_2__N_180[1]), .CK(us_clk), .Q(state[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=14, LSE_LCOL=51, LSE_RCOL=25, LSE_LLINE=76, LSE_RLINE=82 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam state_i1.GSR = "ENABLED";
    FD1P3AX time_high_count_i15 (.D(time_high_count_15__N_183[15]), .SP(us_clk_enable_56), 
            .CK(us_clk), .Q(time_high_count[15])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=51, LSE_RCOL=25, LSE_LLINE=76, LSE_RLINE=82 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i15.GSR = "ENABLED";
    FD1P3AX time_high_count_i14 (.D(time_high_count_15__N_183[14]), .SP(us_clk_enable_56), 
            .CK(us_clk), .Q(time_high_count[14])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=51, LSE_RCOL=25, LSE_LLINE=76, LSE_RLINE=82 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i14.GSR = "ENABLED";
    FD1P3AX time_high_count_i13 (.D(time_high_count_15__N_183[13]), .SP(us_clk_enable_56), 
            .CK(us_clk), .Q(time_high_count[13])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=51, LSE_RCOL=25, LSE_LLINE=76, LSE_RLINE=82 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i13.GSR = "ENABLED";
    FD1P3AX time_high_count_i12 (.D(time_high_count_15__N_183[12]), .SP(us_clk_enable_56), 
            .CK(us_clk), .Q(time_high_count[12])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=51, LSE_RCOL=25, LSE_LLINE=76, LSE_RLINE=82 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i12.GSR = "ENABLED";
    FD1P3AX time_high_count_i11 (.D(time_high_count_15__N_183[11]), .SP(us_clk_enable_56), 
            .CK(us_clk), .Q(time_high_count[11])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=51, LSE_RCOL=25, LSE_LLINE=76, LSE_RLINE=82 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i11.GSR = "ENABLED";
    FD1P3AX time_high_count_i10 (.D(time_high_count_15__N_183[10]), .SP(us_clk_enable_56), 
            .CK(us_clk), .Q(time_high_count[10])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=51, LSE_RCOL=25, LSE_LLINE=76, LSE_RLINE=82 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i10.GSR = "ENABLED";
    FD1P3AX time_high_count_i9 (.D(time_high_count_15__N_183[9]), .SP(us_clk_enable_56), 
            .CK(us_clk), .Q(time_high_count[9])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=51, LSE_RCOL=25, LSE_LLINE=76, LSE_RLINE=82 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i9.GSR = "ENABLED";
    FD1P3AX time_high_count_i8 (.D(time_high_count_15__N_183[8]), .SP(us_clk_enable_56), 
            .CK(us_clk), .Q(time_high_count[8])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=51, LSE_RCOL=25, LSE_LLINE=76, LSE_RLINE=82 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i8.GSR = "ENABLED";
    FD1P3AX time_high_count_i7 (.D(time_high_count_15__N_183[7]), .SP(us_clk_enable_56), 
            .CK(us_clk), .Q(time_high_count[7])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=51, LSE_RCOL=25, LSE_LLINE=76, LSE_RLINE=82 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i7.GSR = "ENABLED";
    FD1P3AX time_high_count_i6 (.D(time_high_count_15__N_183[6]), .SP(us_clk_enable_56), 
            .CK(us_clk), .Q(time_high_count[6])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=51, LSE_RCOL=25, LSE_LLINE=76, LSE_RLINE=82 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i6.GSR = "ENABLED";
    FD1P3AX time_high_count_i5 (.D(time_high_count_15__N_183[5]), .SP(us_clk_enable_56), 
            .CK(us_clk), .Q(time_high_count[5])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=51, LSE_RCOL=25, LSE_LLINE=76, LSE_RLINE=82 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i5.GSR = "ENABLED";
    FD1P3AX time_high_count_i4 (.D(time_high_count_15__N_183[4]), .SP(us_clk_enable_56), 
            .CK(us_clk), .Q(time_high_count[4])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=51, LSE_RCOL=25, LSE_LLINE=76, LSE_RLINE=82 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i4.GSR = "ENABLED";
    FD1P3AX time_high_count_i3 (.D(time_high_count_15__N_183[3]), .SP(us_clk_enable_56), 
            .CK(us_clk), .Q(time_high_count[3])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=51, LSE_RCOL=25, LSE_LLINE=76, LSE_RLINE=82 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i3.GSR = "ENABLED";
    FD1P3AX time_high_count_i2 (.D(time_high_count_15__N_183[2]), .SP(us_clk_enable_58), 
            .CK(us_clk), .Q(time_high_count[2])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=51, LSE_RCOL=25, LSE_LLINE=76, LSE_RLINE=82 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i2.GSR = "ENABLED";
    FD1P3AX time_high_count_i1 (.D(time_high_count_15__N_183[1]), .SP(us_clk_enable_58), 
            .CK(us_clk), .Q(time_high_count[1])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=51, LSE_RCOL=25, LSE_LLINE=76, LSE_RLINE=82 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i1.GSR = "ENABLED";
    LUT4 time_high_count_10__bdd_4_lut_40233 (.A(time_high_count[10]), .B(time_high_count[4]), 
         .C(time_high_count[6]), .D(n52458), .Z(n50712)) /* synthesis lut_function=(A (B+(C (D)))+!A (B (C (D)))) */ ;
    defparam time_high_count_10__bdd_4_lut_40233.init = 16'he888;
    LUT4 time_high_count_10__bdd_2_lut_40234 (.A(time_high_count[10]), .B(time_high_count[4]), 
         .Z(n50713)) /* synthesis lut_function=(A (B)) */ ;
    defparam time_high_count_10__bdd_2_lut_40234.init = 16'h8888;
    LUT4 state_2__N_199_c_1_bdd_4_lut (.A(state_2__N_199_c_1), .B(state[1]), 
         .C(state[0]), .D(pwm_pulse_level_flag), .Z(n51068)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (B+!(C (D))))) */ ;
    defparam state_2__N_199_c_1_bdd_4_lut.init = 16'h1800;
    LUT4 state_2__N_199_c_1_bdd_3_lut (.A(state_2__N_199_c_1), .B(state[1]), 
         .C(state[0]), .Z(n51067)) /* synthesis lut_function=(!(A (B)+!A (B+(C)))) */ ;
    defparam state_2__N_199_c_1_bdd_3_lut.init = 16'h2323;
    LUT4 pwm_pulse_level_flag_I_0_55_1_lut_rep_458 (.A(pwm_pulse_level_flag), 
         .Z(n52394)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[46:74])
    defparam pwm_pulse_level_flag_I_0_55_1_lut_rep_458.init = 16'h5555;
    LUT4 i1_2_lut_2_lut (.A(pwm_pulse_level_flag), .B(state_2__N_199_c_1), 
         .Z(n47221)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[46:74])
    defparam i1_2_lut_2_lut.init = 16'h4444;
    LUT4 i1_3_lut_4_lut (.A(n35569), .B(time_high_count[10]), .C(time_high_count[6]), 
         .D(state[1]), .Z(n3)) /* synthesis lut_function=(A (D)+!A (B (C (D))+!B (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i1_3_lut_4_lut.init = 16'hfb00;
    LUT4 n51112_bdd_3_lut_4_lut (.A(time_high_count[10]), .B(time_high_count[3]), 
         .C(time_high_count[6]), .D(n51111), .Z(n51113)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A ((D)+!C)) */ ;
    defparam n51112_bdd_3_lut_4_lut.init = 16'hfd0d;
    LUT4 time_high_count_10__bdd_2_lut_40237 (.A(time_high_count[10]), .B(time_high_count[3]), 
         .Z(n51110)) /* synthesis lut_function=((B)+!A) */ ;
    defparam time_high_count_10__bdd_2_lut_40237.init = 16'hdddd;
    LUT4 i1_3_lut_4_lut_adj_494 (.A(n35569), .B(time_high_count[10]), .C(time_high_count[7]), 
         .D(state[1]), .Z(n3_adj_5358)) /* synthesis lut_function=(A (D)+!A (B (C (D))+!B (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i1_3_lut_4_lut_adj_494.init = 16'hfb00;
    LUT4 time_high_count_10__bdd_4_lut_40242 (.A(time_high_count[10]), .B(time_high_count[3]), 
         .C(time_high_count[4]), .D(time_high_count[5]), .Z(n51109)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B+!(C (D))))) */ ;
    defparam time_high_count_10__bdd_4_lut_40242.init = 16'h455d;
    LUT4 i1_3_lut_4_lut_adj_495 (.A(n35569), .B(time_high_count[10]), .C(time_high_count[8]), 
         .D(state[1]), .Z(n3_adj_5359)) /* synthesis lut_function=(A (D)+!A (B (C (D))+!B (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i1_3_lut_4_lut_adj_495.init = 16'hfb00;
    LUT4 i1_2_lut_3_lut (.A(n35569), .B(time_high_count[10]), .C(time_high_count[9]), 
         .Z(pwm_pulse_length_us_15__N_208[9])) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i1_2_lut_3_lut.init = 16'hfbfb;
    LUT4 i1_3_lut (.A(n35569), .B(time_high_count[10]), .C(time_high_count[2]), 
         .Z(n152)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i1_3_lut.init = 16'h4040;
    LUT4 i1_2_lut_adj_496 (.A(time_high_count[2]), .B(n35569), .Z(n4)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(57[16:31])
    defparam i1_2_lut_adj_496.init = 16'h2222;
    LUT4 i4_4_lut (.A(n7), .B(time_high_count[12]), .C(time_high_count[13]), 
         .D(time_high_count[14]), .Z(n35569)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i4_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut (.A(time_high_count[11]), .B(time_high_count[15]), .Z(n7)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i39853_3_lut (.A(time_high_count[5]), .B(time_high_count[3]), .C(time_high_count[4]), 
         .Z(n49525)) /* synthesis lut_function=(!(A (B+(C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(57[16:31])
    defparam i39853_3_lut.init = 16'h5757;
    PFUMX i39997 (.BLUT(n50713), .ALUT(n50712), .C0(time_high_count[5]), 
          .Z(n50714));
    PFUMX i40235 (.BLUT(n51110), .ALUT(n51109), .C0(n52458), .Z(n51111));
    LUT4 i21_4_lut (.A(state_2__N_199_c_1), .B(pwm_pulse_level_flag), .C(state[1]), 
         .D(state[0]), .Z(n46791)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A ((D)+!C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(74[13] 161[20])
    defparam i21_4_lut.init = 16'h0a70;
    LUT4 i39917_4_lut (.A(pwm_pulse_level_flag), .B(n48052), .C(state_2__N_199_c_1), 
         .D(state[2]), .Z(us_clk_enable_58)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))))) */ ;
    defparam i39917_4_lut.init = 16'h3337;
    LUT4 i1_2_lut_adj_497 (.A(state[0]), .B(state[1]), .Z(n48052)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_adj_497.init = 16'h2222;
    LUT4 i1_2_lut_adj_498 (.A(state[1]), .B(n35596), .Z(n3_adj_5360)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i1_2_lut_adj_498.init = 16'h8888;
    LUT4 i1_3_lut_adj_499 (.A(n50714), .B(state[1]), .C(n35569), .Z(n3_adj_5361)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i1_3_lut_adj_499.init = 16'hc8c8;
    LUT4 i39451_4_lut (.A(n35569), .B(time_high_count[10]), .C(n62), .D(time_high_count[5]), 
         .Z(pwm_pulse_length_us_15__N_208[5])) /* synthesis lut_function=(!(A+(B (C+!(D))+!B (C (D))))) */ ;
    defparam i39451_4_lut.init = 16'h0511;
    PFUMX i40215 (.BLUT(n51068), .ALUT(n51067), .C0(state[2]), .Z(state_2__N_180[1]));
    LUT4 i39412_3_lut_rep_420 (.A(state[0]), .B(state[1]), .C(state[2]), 
         .Z(us_clk_enable_126)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;
    defparam i39412_3_lut_rep_420.init = 16'hc9c9;
    LUT4 i25776_2_lut (.A(state[2]), .B(state[1]), .Z(n36397)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i25776_2_lut.init = 16'h8888;
    LUT4 i1_4_lut (.A(pwm_pulse_level_flag), .B(state[1]), .C(state_2__N_199_c_1), 
         .D(state[0]), .Z(n46559)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(74[13] 161[20])
    defparam i1_4_lut.init = 16'heccc;
    LUT4 i1_2_lut_4_lut_adj_500 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[15]), .Z(time_high_count_15__N_183[15])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_500.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_501 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[14]), .Z(time_high_count_15__N_183[14])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_501.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_502 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[13]), .Z(time_high_count_15__N_183[13])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_502.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_503 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[12]), .Z(time_high_count_15__N_183[12])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_503.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_504 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[11]), .Z(time_high_count_15__N_183[11])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_504.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_505 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[10]), .Z(time_high_count_15__N_183[10])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_505.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_506 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[9]), .Z(time_high_count_15__N_183[9])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_506.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_507 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[8]), .Z(time_high_count_15__N_183[8])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_507.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_508 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[7]), .Z(time_high_count_15__N_183[7])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_508.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_509 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[6]), .Z(time_high_count_15__N_183[6])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_509.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_510 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[5]), .Z(time_high_count_15__N_183[5])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_510.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_511 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[4]), .Z(time_high_count_15__N_183[4])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_511.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_512 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[3]), .Z(time_high_count_15__N_183[3])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_512.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_513 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[2]), .Z(time_high_count_15__N_183[2])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_513.init = 16'h0400;
    CCU2D add_3747_17 (.A0(n52394), .B0(state_2__N_199_c_1), .C0(time_high_count[15]), 
          .D0(pwm_pulse_level_flag), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43941), .S0(time_high_count_15__N_224[15]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3747_17.INIT0 = 16'hf070;
    defparam add_3747_17.INIT1 = 16'h0000;
    defparam add_3747_17.INJECT1_0 = "NO";
    defparam add_3747_17.INJECT1_1 = "NO";
    CCU2D add_3747_15 (.A0(n52394), .B0(state_2__N_199_c_1), .C0(time_high_count[13]), 
          .D0(pwm_pulse_level_flag), .A1(n52394), .B1(state_2__N_199_c_1), 
          .C1(time_high_count[14]), .D1(pwm_pulse_level_flag), .CIN(n43940), 
          .COUT(n43941), .S0(time_high_count_15__N_224[13]), .S1(time_high_count_15__N_224[14]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3747_15.INIT0 = 16'hf070;
    defparam add_3747_15.INIT1 = 16'hf070;
    defparam add_3747_15.INJECT1_0 = "NO";
    defparam add_3747_15.INJECT1_1 = "NO";
    CCU2D add_3747_13 (.A0(n52394), .B0(state_2__N_199_c_1), .C0(time_high_count[11]), 
          .D0(pwm_pulse_level_flag), .A1(n52394), .B1(state_2__N_199_c_1), 
          .C1(time_high_count[12]), .D1(pwm_pulse_level_flag), .CIN(n43939), 
          .COUT(n43940), .S0(time_high_count_15__N_224[11]), .S1(time_high_count_15__N_224[12]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3747_13.INIT0 = 16'hf070;
    defparam add_3747_13.INIT1 = 16'hf070;
    defparam add_3747_13.INJECT1_0 = "NO";
    defparam add_3747_13.INJECT1_1 = "NO";
    CCU2D add_3747_11 (.A0(n52394), .B0(state_2__N_199_c_1), .C0(time_high_count[9]), 
          .D0(pwm_pulse_level_flag), .A1(n52394), .B1(state_2__N_199_c_1), 
          .C1(time_high_count[10]), .D1(pwm_pulse_level_flag), .CIN(n43938), 
          .COUT(n43939), .S0(time_high_count_15__N_224[9]), .S1(time_high_count_15__N_224[10]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3747_11.INIT0 = 16'hf070;
    defparam add_3747_11.INIT1 = 16'hf070;
    defparam add_3747_11.INJECT1_0 = "NO";
    defparam add_3747_11.INJECT1_1 = "NO";
    CCU2D add_3747_9 (.A0(n52394), .B0(state_2__N_199_c_1), .C0(time_high_count[7]), 
          .D0(pwm_pulse_level_flag), .A1(n52394), .B1(state_2__N_199_c_1), 
          .C1(time_high_count[8]), .D1(pwm_pulse_level_flag), .CIN(n43937), 
          .COUT(n43938), .S0(time_high_count_15__N_224[7]), .S1(time_high_count_15__N_224[8]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3747_9.INIT0 = 16'hf070;
    defparam add_3747_9.INIT1 = 16'hf070;
    defparam add_3747_9.INJECT1_0 = "NO";
    defparam add_3747_9.INJECT1_1 = "NO";
    CCU2D add_3747_7 (.A0(n52394), .B0(state_2__N_199_c_1), .C0(time_high_count[5]), 
          .D0(pwm_pulse_level_flag), .A1(n52394), .B1(state_2__N_199_c_1), 
          .C1(time_high_count[6]), .D1(pwm_pulse_level_flag), .CIN(n43936), 
          .COUT(n43937), .S0(time_high_count_15__N_224[5]), .S1(time_high_count_15__N_224[6]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3747_7.INIT0 = 16'hf070;
    defparam add_3747_7.INIT1 = 16'hf070;
    defparam add_3747_7.INJECT1_0 = "NO";
    defparam add_3747_7.INJECT1_1 = "NO";
    CCU2D add_3747_5 (.A0(n52394), .B0(state_2__N_199_c_1), .C0(time_high_count[3]), 
          .D0(pwm_pulse_level_flag), .A1(n52394), .B1(state_2__N_199_c_1), 
          .C1(time_high_count[4]), .D1(pwm_pulse_level_flag), .CIN(n43935), 
          .COUT(n43936), .S0(time_high_count_15__N_224[3]), .S1(time_high_count_15__N_224[4]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3747_5.INIT0 = 16'hf070;
    defparam add_3747_5.INIT1 = 16'hf070;
    defparam add_3747_5.INJECT1_0 = "NO";
    defparam add_3747_5.INJECT1_1 = "NO";
    CCU2D add_3747_3 (.A0(n52394), .B0(state_2__N_199_c_1), .C0(time_high_count[1]), 
          .D0(pwm_pulse_level_flag), .A1(n52394), .B1(state_2__N_199_c_1), 
          .C1(time_high_count[2]), .D1(pwm_pulse_level_flag), .CIN(n43934), 
          .COUT(n43935), .S0(time_high_count_15__N_224[1]), .S1(time_high_count_15__N_224[2]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3747_3.INIT0 = 16'hf070;
    defparam add_3747_3.INIT1 = 16'hf070;
    defparam add_3747_3.INJECT1_0 = "NO";
    defparam add_3747_3.INJECT1_1 = "NO";
    CCU2D add_3747_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(time_high_count[0]), .B1(n47221), .C1(state_2__N_199_c_1), 
          .D1(pwm_pulse_level_flag), .COUT(n43934), .S1(time_high_count_15__N_224[0]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3747_1.INIT0 = 16'hF000;
    defparam add_3747_1.INIT1 = 16'hd222;
    defparam add_3747_1.INJECT1_0 = "NO";
    defparam add_3747_1.INJECT1_1 = "NO";
    LUT4 i2_3_lut_4_lut (.A(state[1]), .B(state[2]), .C(time_high_count_15__N_224[0]), 
         .D(state[0]), .Z(time_high_count_15__N_183[0])) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i2_3_lut_4_lut.init = 16'h0020;
    LUT4 i20021_2_lut_4_lut_3_lut (.A(state[1]), .B(state[2]), .C(state[0]), 
         .Z(n30688)) /* synthesis lut_function=(A (B)+!A !(B+(C))) */ ;
    defparam i20021_2_lut_4_lut_3_lut.init = 16'h8989;
    LUT4 n51114_bdd_2_lut_3_lut (.A(n51113), .B(state[1]), .C(n35569), 
         .Z(n51115)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam n51114_bdd_2_lut_3_lut.init = 16'h0808;
    PFUMX i24966 (.BLUT(n35593), .ALUT(n35595), .C0(n49525), .Z(n35596));
    LUT4 i2_3_lut_rep_522 (.A(time_high_count[8]), .B(time_high_count[7]), 
         .C(time_high_count[9]), .Z(n52458)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(57[16:31])
    defparam i2_3_lut_rep_522.init = 16'h8080;
    LUT4 i1_2_lut_4_lut_adj_514 (.A(time_high_count[8]), .B(time_high_count[7]), 
         .C(time_high_count[9]), .D(time_high_count[6]), .Z(n80)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(57[16:31])
    defparam i1_2_lut_4_lut_adj_514.init = 16'h8000;
    LUT4 i22_2_lut_4_lut (.A(time_high_count[8]), .B(time_high_count[7]), 
         .C(time_high_count[9]), .D(time_high_count[10]), .Z(n8)) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(57[16:31])
    defparam i22_2_lut_4_lut.init = 16'h7f80;
    FD1P3JX time_high_us_i2 (.D(n3_adj_5360), .SP(us_clk_enable_126), .PD(n30688), 
            .CK(us_clk), .Q(\yaw_pwm_pulse_length_us[2] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=51, LSE_RCOL=25, LSE_LLINE=76, LSE_RLINE=82 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i2.GSR = "ENABLED";
    FD1P3JX time_high_us_i3 (.D(n51115), .SP(us_clk_enable_126), .PD(n30688), 
            .CK(us_clk), .Q(\yaw_pwm_pulse_length_us[3] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=51, LSE_RCOL=25, LSE_LLINE=76, LSE_RLINE=82 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i3.GSR = "ENABLED";
    FD1P3JX time_high_us_i4 (.D(n3_adj_5361), .SP(us_clk_enable_126), .PD(n30688), 
            .CK(us_clk), .Q(\yaw_pwm_pulse_length_us[4] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=51, LSE_RCOL=25, LSE_LLINE=76, LSE_RLINE=82 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i4.GSR = "ENABLED";
    FD1P3IX time_high_us_i5 (.D(pwm_pulse_length_us_15__N_208[5]), .SP(us_clk_enable_126), 
            .CD(n30688), .CK(us_clk), .Q(\yaw_pwm_pulse_length_us[5] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=51, LSE_RCOL=25, LSE_LLINE=76, LSE_RLINE=82 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i5.GSR = "ENABLED";
    FD1P3JX time_high_us_i6 (.D(n3), .SP(us_clk_enable_126), .PD(n30688), 
            .CK(us_clk), .Q(\yaw_pwm_pulse_length_us[6] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=51, LSE_RCOL=25, LSE_LLINE=76, LSE_RLINE=82 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i6.GSR = "ENABLED";
    FD1P3JX time_high_us_i7 (.D(n3_adj_5358), .SP(us_clk_enable_126), .PD(n30688), 
            .CK(us_clk), .Q(\yaw_pwm_pulse_length_us[7] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=51, LSE_RCOL=25, LSE_LLINE=76, LSE_RLINE=82 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i7.GSR = "ENABLED";
    FD1P3JX time_high_us_i8 (.D(n3_adj_5359), .SP(us_clk_enable_126), .PD(n30688), 
            .CK(us_clk), .Q(\yaw_pwm_pulse_length_us[8] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=51, LSE_RCOL=25, LSE_LLINE=76, LSE_RLINE=82 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i8.GSR = "ENABLED";
    FD1P3IX time_high_us_i9 (.D(pwm_pulse_length_us_15__N_208[9]), .SP(us_clk_enable_126), 
            .CD(n30688), .CK(us_clk), .Q(\yaw_pwm_pulse_length_us[9] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=51, LSE_RCOL=25, LSE_LLINE=76, LSE_RLINE=82 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i9.GSR = "ENABLED";
    FD1P3IX pwm_pulse_level_flag_46 (.D(n46559), .SP(us_clk_enable_147), 
            .CD(n36397), .CK(us_clk), .Q(pwm_pulse_level_flag)) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=51, LSE_RCOL=25, LSE_LLINE=76, LSE_RLINE=82 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam pwm_pulse_level_flag_46.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module pwm_to_value
//

module pwm_to_value (yaw_val, us_clk, \yaw_pwm_pulse_length_us[2] , \yaw_pwm_pulse_length_us[5] , 
            \yaw_pwm_pulse_length_us[7] , \yaw_pwm_pulse_length_us[6] , 
            \yaw_pwm_pulse_length_us[8] , \yaw_pwm_pulse_length_us[4] , 
            \yaw_pwm_pulse_length_us[3] , \yaw_pwm_pulse_length_us[9] , 
            n43271, n52456, n51041) /* synthesis syn_module_defined=1 */ ;
    output [7:0]yaw_val;
    input us_clk;
    input \yaw_pwm_pulse_length_us[2] ;
    input \yaw_pwm_pulse_length_us[5] ;
    input \yaw_pwm_pulse_length_us[7] ;
    input \yaw_pwm_pulse_length_us[6] ;
    input \yaw_pwm_pulse_length_us[8] ;
    input \yaw_pwm_pulse_length_us[4] ;
    input \yaw_pwm_pulse_length_us[3] ;
    input \yaw_pwm_pulse_length_us[9] ;
    output n43271;
    output n52456;
    output n51041;
    
    wire us_clk /* synthesis SET_AS_NETWORK=us_clk, is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(221[10:16])
    
    wire n52362;
    wire [15:0]value_out_7__N_154;
    
    wire n52261, n52222;
    
    FD1S3AX adjusted_value_i0 (.D(\yaw_pwm_pulse_length_us[2] ), .CK(us_clk), 
            .Q(yaw_val[0])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=84, LSE_RLINE=89 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i0.GSR = "DISABLED";
    LUT4 i7739_2_lut_3_lut_4_lut (.A(\yaw_pwm_pulse_length_us[5] ), .B(n52362), 
         .C(\yaw_pwm_pulse_length_us[7] ), .D(\yaw_pwm_pulse_length_us[6] ), 
         .Z(value_out_7__N_154[7])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;
    defparam i7739_2_lut_3_lut_4_lut.init = 16'h78f0;
    FD1S3AX adjusted_value_i7 (.D(value_out_7__N_154[9]), .CK(us_clk), .Q(yaw_val[7])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=84, LSE_RLINE=89 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i7.GSR = "DISABLED";
    FD1S3AX adjusted_value_i6 (.D(value_out_7__N_154[8]), .CK(us_clk), .Q(yaw_val[6])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=84, LSE_RLINE=89 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i6.GSR = "DISABLED";
    FD1S3AX adjusted_value_i5 (.D(value_out_7__N_154[7]), .CK(us_clk), .Q(yaw_val[5])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=84, LSE_RLINE=89 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i5.GSR = "DISABLED";
    FD1S3AX adjusted_value_i4 (.D(value_out_7__N_154[6]), .CK(us_clk), .Q(yaw_val[4])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=84, LSE_RLINE=89 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i4.GSR = "DISABLED";
    FD1S3AX adjusted_value_i3 (.D(value_out_7__N_154[5]), .CK(us_clk), .Q(yaw_val[3])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=84, LSE_RLINE=89 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i3.GSR = "DISABLED";
    FD1S3AX adjusted_value_i2 (.D(value_out_7__N_154[4]), .CK(us_clk), .Q(yaw_val[2])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=84, LSE_RLINE=89 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i2.GSR = "DISABLED";
    FD1S3AX adjusted_value_i1 (.D(value_out_7__N_154[3]), .CK(us_clk), .Q(yaw_val[1])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=84, LSE_RLINE=89 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i1.GSR = "DISABLED";
    LUT4 i7746_2_lut_3_lut_4_lut (.A(\yaw_pwm_pulse_length_us[6] ), .B(n52261), 
         .C(\yaw_pwm_pulse_length_us[8] ), .D(\yaw_pwm_pulse_length_us[7] ), 
         .Z(value_out_7__N_154[8])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;
    defparam i7746_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i1_2_lut (.A(\yaw_pwm_pulse_length_us[4] ), .B(\yaw_pwm_pulse_length_us[3] ), 
         .Z(value_out_7__N_154[4])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i1_2_lut.init = 16'h9999;
    LUT4 i7715_1_lut (.A(\yaw_pwm_pulse_length_us[3] ), .Z(value_out_7__N_154[3])) /* synthesis lut_function=(!(A)) */ ;
    defparam i7715_1_lut.init = 16'h5555;
    LUT4 i7753_3_lut_4_lut (.A(\yaw_pwm_pulse_length_us[7] ), .B(n52222), 
         .C(\yaw_pwm_pulse_length_us[8] ), .D(\yaw_pwm_pulse_length_us[9] ), 
         .Z(value_out_7__N_154[9])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;
    defparam i7753_3_lut_4_lut.init = 16'h7f80;
    LUT4 i1_2_lut_2_lut (.A(yaw_val[3]), .B(yaw_val[0]), .Z(n43271)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam i1_2_lut_2_lut.init = 16'hdddd;
    LUT4 i7722_2_lut_rep_426 (.A(\yaw_pwm_pulse_length_us[4] ), .B(\yaw_pwm_pulse_length_us[3] ), 
         .Z(n52362)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i7722_2_lut_rep_426.init = 16'heeee;
    LUT4 i7727_2_lut_rep_325_3_lut (.A(\yaw_pwm_pulse_length_us[4] ), .B(\yaw_pwm_pulse_length_us[3] ), 
         .C(\yaw_pwm_pulse_length_us[5] ), .Z(n52261)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i7727_2_lut_rep_325_3_lut.init = 16'he0e0;
    LUT4 i7725_2_lut_3_lut (.A(\yaw_pwm_pulse_length_us[4] ), .B(\yaw_pwm_pulse_length_us[3] ), 
         .C(\yaw_pwm_pulse_length_us[5] ), .Z(value_out_7__N_154[5])) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B !(C)))) */ ;
    defparam i7725_2_lut_3_lut.init = 16'h1e1e;
    LUT4 i7734_2_lut_rep_286_3_lut_4_lut (.A(\yaw_pwm_pulse_length_us[4] ), 
         .B(\yaw_pwm_pulse_length_us[3] ), .C(\yaw_pwm_pulse_length_us[6] ), 
         .D(\yaw_pwm_pulse_length_us[5] ), .Z(n52222)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;
    defparam i7734_2_lut_rep_286_3_lut_4_lut.init = 16'he000;
    LUT4 i7732_2_lut_3_lut_4_lut (.A(\yaw_pwm_pulse_length_us[4] ), .B(\yaw_pwm_pulse_length_us[3] ), 
         .C(\yaw_pwm_pulse_length_us[6] ), .D(\yaw_pwm_pulse_length_us[5] ), 
         .Z(value_out_7__N_154[6])) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B !(C)))) */ ;
    defparam i7732_2_lut_3_lut_4_lut.init = 16'h1ef0;
    LUT4 i1_2_lut_rep_520 (.A(yaw_val[2]), .B(yaw_val[1]), .Z(n52456)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(77[9:16])
    defparam i1_2_lut_rep_520.init = 16'heeee;
    LUT4 yaw_val_3__bdd_2_lut_40194_3_lut (.A(yaw_val[2]), .B(yaw_val[1]), 
         .C(yaw_val[3]), .Z(n51041)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(77[9:16])
    defparam yaw_val_3__bdd_2_lut_40194_3_lut.init = 16'hefef;
    
endmodule
//
// Verilog Description of module \pwm_reader(DEFAULT_PWM_TIME_HIGH_US=16'b01111101000) 
//

module \pwm_reader(DEFAULT_PWM_TIME_HIGH_US=16'b01111101000)  (state_2__N_84_c_1, 
            GND_net, us_clk, resetn, resetn_derived_2, \i2c_top_debug[1] , 
            n52306, wd_event_active, n52205, n44, n44797, n64, \next_state[0] , 
            n33315, count__auto_time_ms_27__N_1639, n52318, n52142, 
            \i2c_top_debug[5] , byte_rd_left_5__N_1255, \throttle_pwm_pulse_length_us[4] , 
            \throttle_pwm_pulse_length_us[9] , \throttle_pwm_pulse_length_us[8] , 
            \throttle_pwm_pulse_length_us[7] , \throttle_pwm_pulse_length_us[6] , 
            \throttle_pwm_pulse_length_us[5] , \throttle_pwm_pulse_length_us[3] , 
            \throttle_pwm_pulse_length_us[2] ) /* synthesis syn_module_defined=1 */ ;
    input state_2__N_84_c_1;
    input GND_net;
    input us_clk;
    input resetn;
    output resetn_derived_2;
    input \i2c_top_debug[1] ;
    input n52306;
    input wd_event_active;
    output n52205;
    input n44;
    input n44797;
    input n64;
    output \next_state[0] ;
    input n33315;
    output count__auto_time_ms_27__N_1639;
    output n52318;
    input n52142;
    input \i2c_top_debug[5] ;
    output byte_rd_left_5__N_1255;
    output \throttle_pwm_pulse_length_us[4] ;
    output \throttle_pwm_pulse_length_us[9] ;
    output \throttle_pwm_pulse_length_us[8] ;
    output \throttle_pwm_pulse_length_us[7] ;
    output \throttle_pwm_pulse_length_us[6] ;
    output \throttle_pwm_pulse_length_us[5] ;
    output \throttle_pwm_pulse_length_us[3] ;
    output \throttle_pwm_pulse_length_us[2] ;
    
    wire us_clk /* synthesis SET_AS_NETWORK=us_clk, is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(221[10:16])
    wire [2:0]state;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(54[15:20])
    
    wire us_clk_enable_135, n43893, n52307;
    wire [15:0]time_high_count;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(57[16:31])
    
    wire pwm_pulse_level_flag;
    wire [15:0]time_high_count_15__N_109;
    
    wire n43892, n7, n163, n64_c, n43891, n43890, n43889, n43888, 
        n43887, n43886, n47301, n7_adj_5350, n35082, us_clk_enable_94;
    wire [15:0]time_high_count_15__N_68;
    wire [2:0]state_2__N_65;
    
    wire n52305, n47996, n50988, n50989, n52462, n52463, n52034, 
        n48073, us_clk_enable_96, n46753, n52281, n3;
    wire [15:0]pwm_pulse_length_us_15__N_47;
    
    wire n4, us_clk_enable_110, n30785, n51176, n51175, n51177, 
        n125, n52224, n51178, n47993, n36530, n46759, n4_adj_5352, 
        n3_adj_5353, n3_adj_5354, n3_adj_5355, n3_adj_5356;
    
    LUT4 i20_4_lut_3_lut_4_lut (.A(state[1]), .B(state_2__N_84_c_1), .C(state[0]), 
         .D(state[2]), .Z(us_clk_enable_135)) /* synthesis lut_function=(A (B ((D)+!C)+!B (D))+!A !(D)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i20_4_lut_3_lut_4_lut.init = 16'haa5d;
    CCU2D add_3763_17 (.A0(n52307), .B0(state_2__N_84_c_1), .C0(time_high_count[15]), 
          .D0(pwm_pulse_level_flag), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43893), .S0(time_high_count_15__N_109[15]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3763_17.INIT0 = 16'hf070;
    defparam add_3763_17.INIT1 = 16'h0000;
    defparam add_3763_17.INJECT1_0 = "NO";
    defparam add_3763_17.INJECT1_1 = "NO";
    CCU2D add_3763_15 (.A0(n52307), .B0(state_2__N_84_c_1), .C0(time_high_count[13]), 
          .D0(pwm_pulse_level_flag), .A1(n52307), .B1(state_2__N_84_c_1), 
          .C1(time_high_count[14]), .D1(pwm_pulse_level_flag), .CIN(n43892), 
          .COUT(n43893), .S0(time_high_count_15__N_109[13]), .S1(time_high_count_15__N_109[14]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3763_15.INIT0 = 16'hf070;
    defparam add_3763_15.INIT1 = 16'hf070;
    defparam add_3763_15.INJECT1_0 = "NO";
    defparam add_3763_15.INJECT1_1 = "NO";
    PFUMX i45 (.BLUT(n7), .ALUT(n163), .C0(time_high_count[5]), .Z(n64_c));
    CCU2D add_3763_13 (.A0(n52307), .B0(state_2__N_84_c_1), .C0(time_high_count[11]), 
          .D0(pwm_pulse_level_flag), .A1(n52307), .B1(state_2__N_84_c_1), 
          .C1(time_high_count[12]), .D1(pwm_pulse_level_flag), .CIN(n43891), 
          .COUT(n43892), .S0(time_high_count_15__N_109[11]), .S1(time_high_count_15__N_109[12]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3763_13.INIT0 = 16'hf070;
    defparam add_3763_13.INIT1 = 16'hf070;
    defparam add_3763_13.INJECT1_0 = "NO";
    defparam add_3763_13.INJECT1_1 = "NO";
    CCU2D add_3763_11 (.A0(n52307), .B0(state_2__N_84_c_1), .C0(time_high_count[9]), 
          .D0(pwm_pulse_level_flag), .A1(n52307), .B1(state_2__N_84_c_1), 
          .C1(time_high_count[10]), .D1(pwm_pulse_level_flag), .CIN(n43890), 
          .COUT(n43891), .S0(time_high_count_15__N_109[9]), .S1(time_high_count_15__N_109[10]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3763_11.INIT0 = 16'hf070;
    defparam add_3763_11.INIT1 = 16'hf070;
    defparam add_3763_11.INJECT1_0 = "NO";
    defparam add_3763_11.INJECT1_1 = "NO";
    CCU2D add_3763_9 (.A0(n52307), .B0(state_2__N_84_c_1), .C0(time_high_count[7]), 
          .D0(pwm_pulse_level_flag), .A1(n52307), .B1(state_2__N_84_c_1), 
          .C1(time_high_count[8]), .D1(pwm_pulse_level_flag), .CIN(n43889), 
          .COUT(n43890), .S0(time_high_count_15__N_109[7]), .S1(time_high_count_15__N_109[8]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3763_9.INIT0 = 16'hf070;
    defparam add_3763_9.INIT1 = 16'hf070;
    defparam add_3763_9.INJECT1_0 = "NO";
    defparam add_3763_9.INJECT1_1 = "NO";
    CCU2D add_3763_7 (.A0(n52307), .B0(state_2__N_84_c_1), .C0(time_high_count[5]), 
          .D0(pwm_pulse_level_flag), .A1(n52307), .B1(state_2__N_84_c_1), 
          .C1(time_high_count[6]), .D1(pwm_pulse_level_flag), .CIN(n43888), 
          .COUT(n43889), .S0(time_high_count_15__N_109[5]), .S1(time_high_count_15__N_109[6]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3763_7.INIT0 = 16'hf070;
    defparam add_3763_7.INIT1 = 16'hf070;
    defparam add_3763_7.INJECT1_0 = "NO";
    defparam add_3763_7.INJECT1_1 = "NO";
    CCU2D add_3763_5 (.A0(n52307), .B0(state_2__N_84_c_1), .C0(time_high_count[3]), 
          .D0(pwm_pulse_level_flag), .A1(n52307), .B1(state_2__N_84_c_1), 
          .C1(time_high_count[4]), .D1(pwm_pulse_level_flag), .CIN(n43887), 
          .COUT(n43888), .S0(time_high_count_15__N_109[3]), .S1(time_high_count_15__N_109[4]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3763_5.INIT0 = 16'hf070;
    defparam add_3763_5.INIT1 = 16'hf070;
    defparam add_3763_5.INJECT1_0 = "NO";
    defparam add_3763_5.INJECT1_1 = "NO";
    CCU2D add_3763_3 (.A0(n52307), .B0(state_2__N_84_c_1), .C0(time_high_count[1]), 
          .D0(pwm_pulse_level_flag), .A1(n52307), .B1(state_2__N_84_c_1), 
          .C1(time_high_count[2]), .D1(pwm_pulse_level_flag), .CIN(n43886), 
          .COUT(n43887), .S0(time_high_count_15__N_109[1]), .S1(time_high_count_15__N_109[2]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3763_3.INIT0 = 16'hf070;
    defparam add_3763_3.INIT1 = 16'hf070;
    defparam add_3763_3.INJECT1_0 = "NO";
    defparam add_3763_3.INJECT1_1 = "NO";
    CCU2D add_3763_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(time_high_count[0]), .B1(n47301), .C1(state_2__N_84_c_1), 
          .D1(pwm_pulse_level_flag), .COUT(n43886), .S1(time_high_count_15__N_109[0]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3763_1.INIT0 = 16'hF000;
    defparam add_3763_1.INIT1 = 16'hd222;
    defparam add_3763_1.INJECT1_0 = "NO";
    defparam add_3763_1.INJECT1_1 = "NO";
    LUT4 i39655_4_lut (.A(n7_adj_5350), .B(time_high_count[15]), .C(time_high_count[13]), 
         .D(time_high_count[12]), .Z(n35082)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i39655_4_lut.init = 16'h0001;
    LUT4 i2_2_lut (.A(time_high_count[11]), .B(time_high_count[14]), .Z(n7_adj_5350)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i2_2_lut.init = 16'heeee;
    FD1P3AX time_high_count_i0 (.D(time_high_count_15__N_68[0]), .SP(us_clk_enable_94), 
            .CK(us_clk), .Q(time_high_count[0])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=56, LSE_RCOL=25, LSE_LLINE=60, LSE_RLINE=66 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i0.GSR = "ENABLED";
    FD1S3AX state_i0 (.D(state_2__N_65[0]), .CK(us_clk), .Q(state[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=14, LSE_LCOL=56, LSE_RCOL=25, LSE_LLINE=60, LSE_RLINE=66 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam state_i0.GSR = "ENABLED";
    LUT4 i1_3_lut_4_lut (.A(time_high_count[5]), .B(n52305), .C(time_high_count[4]), 
         .D(time_high_count[10]), .Z(n47996)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(57[16:31])
    defparam i1_3_lut_4_lut.init = 16'h8880;
    LUT4 state_2__N_84_c_1_bdd_3_lut (.A(state_2__N_84_c_1), .B(state[1]), 
         .C(state[0]), .Z(n50988)) /* synthesis lut_function=(!(A (B)+!A (B+(C)))) */ ;
    defparam state_2__N_84_c_1_bdd_3_lut.init = 16'h2323;
    LUT4 state_2__N_84_c_1_bdd_4_lut (.A(state_2__N_84_c_1), .B(state[1]), 
         .C(state[0]), .D(pwm_pulse_level_flag), .Z(n50989)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (B+!(C (D))))) */ ;
    defparam state_2__N_84_c_1_bdd_4_lut.init = 16'h1800;
    LUT4 i1_2_lut_rep_526 (.A(time_high_count[6]), .B(time_high_count[9]), 
         .Z(n52462)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(57[16:31])
    defparam i1_2_lut_rep_526.init = 16'h8888;
    LUT4 time_high_count_4__bdd_4_lut (.A(time_high_count[4]), .B(n52463), 
         .C(time_high_count[3]), .D(time_high_count[10]), .Z(n52034)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B ((D)+!C)+!B !(D)))) */ ;
    defparam time_high_count_4__bdd_4_lut.init = 16'h33c8;
    LUT4 pwm_pulse_level_flag_I_0_55_1_lut_rep_371 (.A(pwm_pulse_level_flag), 
         .Z(n52307)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[46:74])
    defparam pwm_pulse_level_flag_I_0_55_1_lut_rep_371.init = 16'h5555;
    LUT4 i1_2_lut_2_lut (.A(pwm_pulse_level_flag), .B(state_2__N_84_c_1), 
         .Z(n47301)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[46:74])
    defparam i1_2_lut_2_lut.init = 16'h4444;
    LUT4 resetn_I_0_743_1_lut_rep_381 (.A(resetn), .Z(resetn_derived_2)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(242[12:19])
    defparam resetn_I_0_743_1_lut_rep_381.init = 16'h5555;
    LUT4 i39877_2_lut_rep_269_3_lut_4_lut_4_lut (.A(resetn), .B(\i2c_top_debug[1] ), 
         .C(n52306), .D(wd_event_active), .Z(n52205)) /* synthesis lut_function=(!((B (D)+!B ((D)+!C))+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(242[12:19])
    defparam i39877_2_lut_rep_269_3_lut_4_lut_4_lut.init = 16'h00a8;
    LUT4 i1_4_lut_4_lut (.A(resetn), .B(n44), .C(n44797), .D(n64), .Z(\next_state[0] )) /* synthesis lut_function=((B (C)+!B !(D))+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(242[12:19])
    defparam i1_4_lut_4_lut.init = 16'hd5f7;
    LUT4 i1_2_lut_2_lut_adj_469 (.A(resetn), .B(n33315), .Z(count__auto_time_ms_27__N_1639)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(242[12:19])
    defparam i1_2_lut_2_lut_adj_469.init = 16'hdddd;
    LUT4 i11353_2_lut_rep_382 (.A(resetn), .B(wd_event_active), .Z(n52318)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(242[12:19])
    defparam i11353_2_lut_rep_382.init = 16'hdddd;
    LUT4 i39632_4_lut_4_lut (.A(resetn), .B(wd_event_active), .C(n52142), 
         .D(\i2c_top_debug[5] ), .Z(byte_rd_left_5__N_1255)) /* synthesis lut_function=(!(A (B+(C+(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(242[12:19])
    defparam i39632_4_lut_4_lut.init = 16'h5557;
    LUT4 i39676_4_lut (.A(pwm_pulse_level_flag), .B(n48073), .C(state_2__N_84_c_1), 
         .D(state[2]), .Z(us_clk_enable_96)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))))) */ ;
    defparam i39676_4_lut.init = 16'h3337;
    LUT4 i21_4_lut (.A(state_2__N_84_c_1), .B(pwm_pulse_level_flag), .C(state[1]), 
         .D(state[0]), .Z(n46753)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A ((D)+!C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(74[13] 161[20])
    defparam i21_4_lut.init = 16'h0a70;
    LUT4 i1_4_lut (.A(n47996), .B(n52281), .C(n35082), .D(n3), .Z(pwm_pulse_length_us_15__N_47[4])) /* synthesis lut_function=(!(A (B)+!A (B+!((D)+!C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i1_4_lut.init = 16'h3323;
    LUT4 i1_2_lut (.A(time_high_count[10]), .B(time_high_count[4]), .Z(n3)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_4_lut (.A(state[2]), .B(state[1]), .C(state[0]), .D(time_high_count_15__N_109[0]), 
         .Z(time_high_count_15__N_68[0])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_470 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_109[1]), .Z(time_high_count_15__N_68[1])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_470.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_471 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_109[2]), .Z(time_high_count_15__N_68[2])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_471.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_472 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_109[3]), .Z(time_high_count_15__N_68[3])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_472.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_473 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_109[4]), .Z(time_high_count_15__N_68[4])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_473.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_474 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_109[5]), .Z(time_high_count_15__N_68[5])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_474.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_475 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_109[6]), .Z(time_high_count_15__N_68[6])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_475.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_476 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_109[7]), .Z(time_high_count_15__N_68[7])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_476.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_477 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_109[8]), .Z(time_high_count_15__N_68[8])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_477.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_478 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_109[9]), .Z(time_high_count_15__N_68[9])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_478.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_479 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_109[10]), .Z(time_high_count_15__N_68[10])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_479.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_480 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_109[11]), .Z(time_high_count_15__N_68[11])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_480.init = 16'h0400;
    LUT4 i1_2_lut_adj_481 (.A(state[0]), .B(state[1]), .Z(n48073)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_adj_481.init = 16'h2222;
    LUT4 i1_2_lut_4_lut_adj_482 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_109[12]), .Z(time_high_count_15__N_68[12])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_482.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_483 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_109[13]), .Z(time_high_count_15__N_68[13])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_483.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_484 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_109[14]), .Z(time_high_count_15__N_68[14])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_484.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_485 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_109[15]), .Z(time_high_count_15__N_68[15])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_485.init = 16'h0400;
    LUT4 i2_4_lut (.A(state[0]), .B(state_2__N_84_c_1), .C(state[1]), 
         .D(n4), .Z(us_clk_enable_94)) /* synthesis lut_function=((B (C)+!B (C+!(D)))+!A) */ ;
    defparam i2_4_lut.init = 16'hf5f7;
    LUT4 i1_2_lut_adj_486 (.A(state[2]), .B(pwm_pulse_level_flag), .Z(n4)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_486.init = 16'heeee;
    LUT4 i39414_3_lut_rep_481 (.A(state[0]), .B(state[1]), .C(state[2]), 
         .Z(us_clk_enable_110)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;
    defparam i39414_3_lut_rep_481.init = 16'hc9c9;
    LUT4 i20114_2_lut_3_lut_3_lut_3_lut (.A(state[0]), .B(state[1]), .C(state[2]), 
         .Z(n30785)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B !(C))) */ ;
    defparam i20114_2_lut_3_lut_3_lut_3_lut.init = 16'hc1c1;
    PFUMX i40272 (.BLUT(n51176), .ALUT(n51175), .C0(n52305), .Z(n51177));
    LUT4 n149_bdd_2_lut_40287 (.A(time_high_count[3]), .B(time_high_count[10]), 
         .Z(n51176)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam n149_bdd_2_lut_40287.init = 16'hbbbb;
    LUT4 n149_bdd_4_lut_40286 (.A(time_high_count[3]), .B(time_high_count[5]), 
         .C(time_high_count[4]), .D(time_high_count[10]), .Z(n51175)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)))+!A (B (C+(D))+!B (D)))) */ ;
    defparam n149_bdd_4_lut_40286.init = 16'h02bf;
    LUT4 i1_2_lut_3_lut (.A(time_high_count[6]), .B(time_high_count[9]), 
         .C(time_high_count[4]), .Z(n125)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(57[16:31])
    defparam i1_2_lut_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_288 (.A(state[1]), .B(n35082), .Z(n52224)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_288.init = 16'h8888;
    LUT4 gnd_bdd_2_lut_40294_3_lut (.A(state[1]), .B(n35082), .C(n51177), 
         .Z(n51178)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam gnd_bdd_2_lut_40294_3_lut.init = 16'h8080;
    LUT4 i1_4_lut_adj_487 (.A(time_high_count[5]), .B(n52224), .C(time_high_count[10]), 
         .D(n52305), .Z(n47993)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A ((C)+!B))) */ ;
    defparam i1_4_lut_adj_487.init = 16'h0c8c;
    LUT4 state_2__N_84_c_1_bdd_4_lut_40162 (.A(state_2__N_84_c_1), .B(state[2]), 
         .C(state[0]), .D(state[1]), .Z(state_2__N_65[0])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B ((D)+!C)))) */ ;
    defparam state_2__N_84_c_1_bdd_4_lut_40162.init = 16'h3173;
    FD1P3AX time_high_count_i1 (.D(time_high_count_15__N_68[1]), .SP(us_clk_enable_94), 
            .CK(us_clk), .Q(time_high_count[1])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=56, LSE_RCOL=25, LSE_LLINE=60, LSE_RLINE=66 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i1.GSR = "ENABLED";
    FD1P3AX time_high_count_i2 (.D(time_high_count_15__N_68[2]), .SP(us_clk_enable_94), 
            .CK(us_clk), .Q(time_high_count[2])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=56, LSE_RCOL=25, LSE_LLINE=60, LSE_RLINE=66 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i2.GSR = "ENABLED";
    FD1P3AX time_high_count_i3 (.D(time_high_count_15__N_68[3]), .SP(us_clk_enable_94), 
            .CK(us_clk), .Q(time_high_count[3])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=56, LSE_RCOL=25, LSE_LLINE=60, LSE_RLINE=66 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i3.GSR = "ENABLED";
    FD1P3AX time_high_count_i4 (.D(time_high_count_15__N_68[4]), .SP(us_clk_enable_94), 
            .CK(us_clk), .Q(time_high_count[4])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=56, LSE_RCOL=25, LSE_LLINE=60, LSE_RLINE=66 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i4.GSR = "ENABLED";
    FD1P3AX time_high_count_i5 (.D(time_high_count_15__N_68[5]), .SP(us_clk_enable_94), 
            .CK(us_clk), .Q(time_high_count[5])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=56, LSE_RCOL=25, LSE_LLINE=60, LSE_RLINE=66 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i5.GSR = "ENABLED";
    FD1P3AX time_high_count_i6 (.D(time_high_count_15__N_68[6]), .SP(us_clk_enable_94), 
            .CK(us_clk), .Q(time_high_count[6])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=56, LSE_RCOL=25, LSE_LLINE=60, LSE_RLINE=66 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i6.GSR = "ENABLED";
    FD1P3AX time_high_count_i7 (.D(time_high_count_15__N_68[7]), .SP(us_clk_enable_94), 
            .CK(us_clk), .Q(time_high_count[7])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=56, LSE_RCOL=25, LSE_LLINE=60, LSE_RLINE=66 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i7.GSR = "ENABLED";
    FD1P3AX time_high_count_i8 (.D(time_high_count_15__N_68[8]), .SP(us_clk_enable_94), 
            .CK(us_clk), .Q(time_high_count[8])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=56, LSE_RCOL=25, LSE_LLINE=60, LSE_RLINE=66 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i8.GSR = "ENABLED";
    FD1P3AX time_high_count_i9 (.D(time_high_count_15__N_68[9]), .SP(us_clk_enable_94), 
            .CK(us_clk), .Q(time_high_count[9])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=56, LSE_RCOL=25, LSE_LLINE=60, LSE_RLINE=66 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i9.GSR = "ENABLED";
    FD1P3AX time_high_count_i10 (.D(time_high_count_15__N_68[10]), .SP(us_clk_enable_94), 
            .CK(us_clk), .Q(time_high_count[10])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=56, LSE_RCOL=25, LSE_LLINE=60, LSE_RLINE=66 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i10.GSR = "ENABLED";
    FD1P3AX time_high_count_i11 (.D(time_high_count_15__N_68[11]), .SP(us_clk_enable_94), 
            .CK(us_clk), .Q(time_high_count[11])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=56, LSE_RCOL=25, LSE_LLINE=60, LSE_RLINE=66 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i11.GSR = "ENABLED";
    FD1P3AX time_high_count_i12 (.D(time_high_count_15__N_68[12]), .SP(us_clk_enable_94), 
            .CK(us_clk), .Q(time_high_count[12])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=56, LSE_RCOL=25, LSE_LLINE=60, LSE_RLINE=66 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i12.GSR = "ENABLED";
    FD1P3AX time_high_count_i13 (.D(time_high_count_15__N_68[13]), .SP(us_clk_enable_94), 
            .CK(us_clk), .Q(time_high_count[13])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=56, LSE_RCOL=25, LSE_LLINE=60, LSE_RLINE=66 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i13.GSR = "ENABLED";
    FD1P3AX time_high_count_i14 (.D(time_high_count_15__N_68[14]), .SP(us_clk_enable_96), 
            .CK(us_clk), .Q(time_high_count[14])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=56, LSE_RCOL=25, LSE_LLINE=60, LSE_RLINE=66 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i14.GSR = "ENABLED";
    FD1P3AX time_high_count_i15 (.D(time_high_count_15__N_68[15]), .SP(us_clk_enable_96), 
            .CK(us_clk), .Q(time_high_count[15])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=56, LSE_RCOL=25, LSE_LLINE=60, LSE_RLINE=66 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i15.GSR = "ENABLED";
    FD1S3AX state_i1 (.D(state_2__N_65[1]), .CK(us_clk), .Q(state[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=14, LSE_LCOL=56, LSE_RCOL=25, LSE_LLINE=60, LSE_RLINE=66 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam state_i1.GSR = "ENABLED";
    FD1S3IX state_i2 (.D(n46753), .CK(us_clk), .CD(state[2]), .Q(state[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=14, LSE_LCOL=56, LSE_RCOL=25, LSE_LLINE=60, LSE_RLINE=66 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam state_i2.GSR = "ENABLED";
    FD1P3AX time_high_us_i4 (.D(pwm_pulse_length_us_15__N_47[4]), .SP(us_clk_enable_110), 
            .CK(us_clk), .Q(\throttle_pwm_pulse_length_us[4] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=56, LSE_RCOL=25, LSE_LLINE=60, LSE_RLINE=66 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i4.GSR = "ENABLED";
    LUT4 i25908_2_lut (.A(state[2]), .B(state[1]), .Z(n36530)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i25908_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_488 (.A(pwm_pulse_level_flag), .B(state[1]), .C(state_2__N_84_c_1), 
         .D(state[0]), .Z(n46759)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(74[13] 161[20])
    defparam i1_4_lut_adj_488.init = 16'heccc;
    PFUMX i40163 (.BLUT(n50989), .ALUT(n50988), .C0(state[2]), .Z(state_2__N_65[1]));
    LUT4 i155_2_lut_rep_345_2_lut (.A(state[1]), .B(state[2]), .Z(n52281)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i155_2_lut_rep_345_2_lut.init = 16'hdddd;
    LUT4 i2_3_lut_4_lut_4_lut (.A(state[1]), .B(time_high_count[2]), .C(n64_c), 
         .D(state[2]), .Z(pwm_pulse_length_us_15__N_47[2])) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i2_3_lut_4_lut_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_rep_527 (.A(time_high_count[7]), .B(time_high_count[8]), 
         .Z(n52463)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i1_2_lut_rep_527.init = 16'h8888;
    LUT4 i1_2_lut_rep_369_3_lut_4_lut (.A(time_high_count[7]), .B(time_high_count[8]), 
         .C(time_high_count[9]), .D(time_high_count[6]), .Z(n52305)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i1_2_lut_rep_369_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_adj_489 (.A(time_high_count[7]), .B(time_high_count[8]), 
         .C(time_high_count[10]), .Z(n4_adj_5352)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i1_2_lut_3_lut_adj_489.init = 16'h7070;
    LUT4 i154_4_lut_4_lut (.A(time_high_count[10]), .B(n35082), .C(n52034), 
         .D(n52462), .Z(n163)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i154_4_lut_4_lut.init = 16'hc088;
    LUT4 i1_3_lut_4_lut_adj_490 (.A(time_high_count[10]), .B(n35082), .C(time_high_count[9]), 
         .D(state[1]), .Z(n3_adj_5353)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (D)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i1_3_lut_4_lut_adj_490.init = 16'hf700;
    LUT4 i41_4_lut_4_lut (.A(time_high_count[10]), .B(n35082), .C(n4_adj_5352), 
         .D(n125), .Z(n7)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i41_4_lut_4_lut.init = 16'hc088;
    LUT4 i1_3_lut_4_lut_adj_491 (.A(time_high_count[10]), .B(n35082), .C(time_high_count[8]), 
         .D(state[1]), .Z(n3_adj_5354)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (D)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i1_3_lut_4_lut_adj_491.init = 16'hf700;
    LUT4 i1_3_lut_4_lut_adj_492 (.A(time_high_count[10]), .B(n35082), .C(time_high_count[7]), 
         .D(state[1]), .Z(n3_adj_5355)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (D)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i1_3_lut_4_lut_adj_492.init = 16'hf700;
    FD1P3JX time_high_us_i9 (.D(n3_adj_5353), .SP(us_clk_enable_110), .PD(n30785), 
            .CK(us_clk), .Q(\throttle_pwm_pulse_length_us[9] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=56, LSE_RCOL=25, LSE_LLINE=60, LSE_RLINE=66 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i9.GSR = "ENABLED";
    FD1P3JX time_high_us_i8 (.D(n3_adj_5354), .SP(us_clk_enable_110), .PD(n30785), 
            .CK(us_clk), .Q(\throttle_pwm_pulse_length_us[8] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=56, LSE_RCOL=25, LSE_LLINE=60, LSE_RLINE=66 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i8.GSR = "ENABLED";
    FD1P3JX time_high_us_i7 (.D(n3_adj_5355), .SP(us_clk_enable_110), .PD(n30785), 
            .CK(us_clk), .Q(\throttle_pwm_pulse_length_us[7] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=56, LSE_RCOL=25, LSE_LLINE=60, LSE_RLINE=66 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i7.GSR = "ENABLED";
    FD1P3JX time_high_us_i6 (.D(n3_adj_5356), .SP(us_clk_enable_110), .PD(n30785), 
            .CK(us_clk), .Q(\throttle_pwm_pulse_length_us[6] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=56, LSE_RCOL=25, LSE_LLINE=60, LSE_RLINE=66 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i6.GSR = "ENABLED";
    FD1P3JX time_high_us_i5 (.D(n47993), .SP(us_clk_enable_110), .PD(n30785), 
            .CK(us_clk), .Q(\throttle_pwm_pulse_length_us[5] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=56, LSE_RCOL=25, LSE_LLINE=60, LSE_RLINE=66 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i5.GSR = "ENABLED";
    FD1P3JX time_high_us_i3 (.D(n51178), .SP(us_clk_enable_110), .PD(n30785), 
            .CK(us_clk), .Q(\throttle_pwm_pulse_length_us[3] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=56, LSE_RCOL=25, LSE_LLINE=60, LSE_RLINE=66 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i3.GSR = "ENABLED";
    FD1P3AX time_high_us_i2 (.D(pwm_pulse_length_us_15__N_47[2]), .SP(us_clk_enable_110), 
            .CK(us_clk), .Q(\throttle_pwm_pulse_length_us[2] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=56, LSE_RCOL=25, LSE_LLINE=60, LSE_RLINE=66 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i2.GSR = "ENABLED";
    FD1P3IX pwm_pulse_level_flag_46 (.D(n46759), .SP(us_clk_enable_135), 
            .CD(n36530), .CK(us_clk), .Q(pwm_pulse_level_flag)) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=56, LSE_RCOL=25, LSE_LLINE=60, LSE_RLINE=66 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam pwm_pulse_level_flag_46.GSR = "ENABLED";
    LUT4 i1_3_lut_4_lut_adj_493 (.A(time_high_count[10]), .B(n35082), .C(time_high_count[6]), 
         .D(state[1]), .Z(n3_adj_5356)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (D)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i1_3_lut_4_lut_adj_493.init = 16'hf700;
    
endmodule
//
// Verilog Description of module pwm_to_value_U0
//

module pwm_to_value_U0 (throttle_val, us_clk, \throttle_pwm_pulse_length_us[2] , 
            \throttle_pwm_pulse_length_us[5] , \throttle_pwm_pulse_length_us[7] , 
            \throttle_pwm_pulse_length_us[6] , \throttle_pwm_pulse_length_us[8] , 
            n52441, n51044, \throttle_pwm_pulse_length_us[9] , \throttle_pwm_pulse_length_us[4] , 
            \throttle_pwm_pulse_length_us[3] , n52429) /* synthesis syn_module_defined=1 */ ;
    output [7:0]throttle_val;
    input us_clk;
    input \throttle_pwm_pulse_length_us[2] ;
    input \throttle_pwm_pulse_length_us[5] ;
    input \throttle_pwm_pulse_length_us[7] ;
    input \throttle_pwm_pulse_length_us[6] ;
    input \throttle_pwm_pulse_length_us[8] ;
    output n52441;
    output n51044;
    input \throttle_pwm_pulse_length_us[9] ;
    input \throttle_pwm_pulse_length_us[4] ;
    input \throttle_pwm_pulse_length_us[3] ;
    output n52429;
    
    wire us_clk /* synthesis SET_AS_NETWORK=us_clk, is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(221[10:16])
    
    wire n52355;
    wire [15:0]value_out_7__N_154;
    
    wire n52260, n52221;
    
    FD1S3AX adjusted_value_i0 (.D(\throttle_pwm_pulse_length_us[2] ), .CK(us_clk), 
            .Q(throttle_val[0])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=68, LSE_RLINE=73 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i0.GSR = "DISABLED";
    LUT4 i7557_2_lut_3_lut_4_lut (.A(\throttle_pwm_pulse_length_us[5] ), .B(n52355), 
         .C(\throttle_pwm_pulse_length_us[7] ), .D(\throttle_pwm_pulse_length_us[6] ), 
         .Z(value_out_7__N_154[7])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;
    defparam i7557_2_lut_3_lut_4_lut.init = 16'h78f0;
    FD1S3AX adjusted_value_i7 (.D(value_out_7__N_154[9]), .CK(us_clk), .Q(throttle_val[7])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=68, LSE_RLINE=73 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i7.GSR = "DISABLED";
    FD1S3AX adjusted_value_i6 (.D(value_out_7__N_154[8]), .CK(us_clk), .Q(throttle_val[6])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=68, LSE_RLINE=73 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i6.GSR = "DISABLED";
    FD1S3AX adjusted_value_i5 (.D(value_out_7__N_154[7]), .CK(us_clk), .Q(throttle_val[5])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=68, LSE_RLINE=73 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i5.GSR = "DISABLED";
    FD1S3AX adjusted_value_i4 (.D(value_out_7__N_154[6]), .CK(us_clk), .Q(throttle_val[4])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=68, LSE_RLINE=73 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i4.GSR = "DISABLED";
    FD1S3AX adjusted_value_i3 (.D(value_out_7__N_154[5]), .CK(us_clk), .Q(throttle_val[3])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=68, LSE_RLINE=73 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i3.GSR = "DISABLED";
    FD1S3AX adjusted_value_i2 (.D(value_out_7__N_154[4]), .CK(us_clk), .Q(throttle_val[2])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=68, LSE_RLINE=73 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i2.GSR = "DISABLED";
    FD1S3AX adjusted_value_i1 (.D(value_out_7__N_154[3]), .CK(us_clk), .Q(throttle_val[1])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=68, LSE_RLINE=73 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i1.GSR = "DISABLED";
    LUT4 i7564_2_lut_3_lut_4_lut (.A(\throttle_pwm_pulse_length_us[6] ), .B(n52260), 
         .C(\throttle_pwm_pulse_length_us[8] ), .D(\throttle_pwm_pulse_length_us[7] ), 
         .Z(value_out_7__N_154[8])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;
    defparam i7564_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i1_2_lut_rep_505 (.A(throttle_val[1]), .B(throttle_val[2]), .Z(n52441)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(76[9:21])
    defparam i1_2_lut_rep_505.init = 16'heeee;
    LUT4 n48138_bdd_2_lut_40197_3_lut (.A(throttle_val[1]), .B(throttle_val[2]), 
         .C(throttle_val[3]), .Z(n51044)) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(76[9:21])
    defparam n48138_bdd_2_lut_40197_3_lut.init = 16'hefef;
    LUT4 i7571_3_lut_4_lut (.A(\throttle_pwm_pulse_length_us[7] ), .B(n52221), 
         .C(\throttle_pwm_pulse_length_us[8] ), .D(\throttle_pwm_pulse_length_us[9] ), 
         .Z(value_out_7__N_154[9])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;
    defparam i7571_3_lut_4_lut.init = 16'h7f80;
    LUT4 i1_2_lut (.A(\throttle_pwm_pulse_length_us[4] ), .B(\throttle_pwm_pulse_length_us[3] ), 
         .Z(value_out_7__N_154[4])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i1_2_lut.init = 16'h9999;
    LUT4 i7533_1_lut (.A(\throttle_pwm_pulse_length_us[3] ), .Z(value_out_7__N_154[3])) /* synthesis lut_function=(!(A)) */ ;
    defparam i7533_1_lut.init = 16'h5555;
    LUT4 i7540_2_lut_rep_419 (.A(\throttle_pwm_pulse_length_us[4] ), .B(\throttle_pwm_pulse_length_us[3] ), 
         .Z(n52355)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i7540_2_lut_rep_419.init = 16'heeee;
    LUT4 i7545_2_lut_rep_324_3_lut (.A(\throttle_pwm_pulse_length_us[4] ), 
         .B(\throttle_pwm_pulse_length_us[3] ), .C(\throttle_pwm_pulse_length_us[5] ), 
         .Z(n52260)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i7545_2_lut_rep_324_3_lut.init = 16'he0e0;
    LUT4 i7543_2_lut_3_lut (.A(\throttle_pwm_pulse_length_us[4] ), .B(\throttle_pwm_pulse_length_us[3] ), 
         .C(\throttle_pwm_pulse_length_us[5] ), .Z(value_out_7__N_154[5])) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B !(C)))) */ ;
    defparam i7543_2_lut_3_lut.init = 16'h1e1e;
    LUT4 i7552_2_lut_rep_285_3_lut_4_lut (.A(\throttle_pwm_pulse_length_us[4] ), 
         .B(\throttle_pwm_pulse_length_us[3] ), .C(\throttle_pwm_pulse_length_us[6] ), 
         .D(\throttle_pwm_pulse_length_us[5] ), .Z(n52221)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;
    defparam i7552_2_lut_rep_285_3_lut_4_lut.init = 16'he000;
    LUT4 i7550_2_lut_3_lut_4_lut (.A(\throttle_pwm_pulse_length_us[4] ), .B(\throttle_pwm_pulse_length_us[3] ), 
         .C(\throttle_pwm_pulse_length_us[6] ), .D(\throttle_pwm_pulse_length_us[5] ), 
         .Z(value_out_7__N_154[6])) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B !(C)))) */ ;
    defparam i7550_2_lut_3_lut_4_lut.init = 16'h1ef0;
    LUT4 i1_2_lut_rep_493 (.A(throttle_val[3]), .B(throttle_val[0]), .Z(n52429)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam i1_2_lut_rep_493.init = 16'hdddd;
    
endmodule
//
// Verilog Description of module pwm_to_value_U1
//

module pwm_to_value_U1 (\swa_swb_pwm_pulse_length_us[5] , \swa_swb_pwm_pulse_length_us[7] , 
            \swa_swb_pwm_pulse_length_us[6] , swa_swb_val, us_clk, \swa_swb_pwm_pulse_length_us[2] , 
            \swa_swb_pwm_pulse_length_us[8] , \swa_swb_pwm_pulse_length_us[9] , 
            \swa_swb_pwm_pulse_length_us[4] , \swa_swb_pwm_pulse_length_us[3] ) /* synthesis syn_module_defined=1 */ ;
    input \swa_swb_pwm_pulse_length_us[5] ;
    input \swa_swb_pwm_pulse_length_us[7] ;
    input \swa_swb_pwm_pulse_length_us[6] ;
    output [7:0]swa_swb_val;
    input us_clk;
    input \swa_swb_pwm_pulse_length_us[2] ;
    input \swa_swb_pwm_pulse_length_us[8] ;
    input \swa_swb_pwm_pulse_length_us[9] ;
    input \swa_swb_pwm_pulse_length_us[4] ;
    input \swa_swb_pwm_pulse_length_us[3] ;
    
    wire us_clk /* synthesis SET_AS_NETWORK=us_clk, is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(221[10:16])
    
    wire n52327;
    wire [15:0]value_out_7__N_154;
    
    wire n52253, n52215;
    
    LUT4 i7506_2_lut_3_lut_4_lut (.A(\swa_swb_pwm_pulse_length_us[5] ), .B(n52327), 
         .C(\swa_swb_pwm_pulse_length_us[7] ), .D(\swa_swb_pwm_pulse_length_us[6] ), 
         .Z(value_out_7__N_154[7])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;
    defparam i7506_2_lut_3_lut_4_lut.init = 16'h78f0;
    FD1S3AX adjusted_value_i0 (.D(\swa_swb_pwm_pulse_length_us[2] ), .CK(us_clk), 
            .Q(swa_swb_val[0])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=167, LSE_RLINE=172 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i0.GSR = "DISABLED";
    LUT4 i7513_2_lut_3_lut_4_lut (.A(\swa_swb_pwm_pulse_length_us[6] ), .B(n52253), 
         .C(\swa_swb_pwm_pulse_length_us[8] ), .D(\swa_swb_pwm_pulse_length_us[7] ), 
         .Z(value_out_7__N_154[8])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;
    defparam i7513_2_lut_3_lut_4_lut.init = 16'h78f0;
    FD1S3AX adjusted_value_i7 (.D(value_out_7__N_154[9]), .CK(us_clk), .Q(swa_swb_val[7])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=167, LSE_RLINE=172 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i7.GSR = "DISABLED";
    FD1S3AX adjusted_value_i6 (.D(value_out_7__N_154[8]), .CK(us_clk), .Q(swa_swb_val[6])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=167, LSE_RLINE=172 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i6.GSR = "DISABLED";
    FD1S3AX adjusted_value_i5 (.D(value_out_7__N_154[7]), .CK(us_clk), .Q(swa_swb_val[5])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=167, LSE_RLINE=172 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i5.GSR = "DISABLED";
    FD1S3AX adjusted_value_i4 (.D(value_out_7__N_154[6]), .CK(us_clk), .Q(swa_swb_val[4])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=167, LSE_RLINE=172 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i4.GSR = "DISABLED";
    LUT4 i7520_3_lut_4_lut (.A(\swa_swb_pwm_pulse_length_us[7] ), .B(n52215), 
         .C(\swa_swb_pwm_pulse_length_us[8] ), .D(\swa_swb_pwm_pulse_length_us[9] ), 
         .Z(value_out_7__N_154[9])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;
    defparam i7520_3_lut_4_lut.init = 16'h7f80;
    FD1S3AX adjusted_value_i3 (.D(value_out_7__N_154[5]), .CK(us_clk), .Q(swa_swb_val[3])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=167, LSE_RLINE=172 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i3.GSR = "DISABLED";
    FD1S3AX adjusted_value_i2 (.D(value_out_7__N_154[4]), .CK(us_clk), .Q(swa_swb_val[2])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=167, LSE_RLINE=172 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i2.GSR = "DISABLED";
    FD1S3AX adjusted_value_i1 (.D(value_out_7__N_154[3]), .CK(us_clk), .Q(swa_swb_val[1])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=167, LSE_RLINE=172 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i1.GSR = "DISABLED";
    LUT4 i7489_2_lut_rep_391 (.A(\swa_swb_pwm_pulse_length_us[4] ), .B(\swa_swb_pwm_pulse_length_us[3] ), 
         .Z(n52327)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i7489_2_lut_rep_391.init = 16'heeee;
    LUT4 i7494_2_lut_rep_317_3_lut (.A(\swa_swb_pwm_pulse_length_us[4] ), 
         .B(\swa_swb_pwm_pulse_length_us[3] ), .C(\swa_swb_pwm_pulse_length_us[5] ), 
         .Z(n52253)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i7494_2_lut_rep_317_3_lut.init = 16'he0e0;
    LUT4 i7492_2_lut_3_lut (.A(\swa_swb_pwm_pulse_length_us[4] ), .B(\swa_swb_pwm_pulse_length_us[3] ), 
         .C(\swa_swb_pwm_pulse_length_us[5] ), .Z(value_out_7__N_154[5])) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B !(C)))) */ ;
    defparam i7492_2_lut_3_lut.init = 16'h1e1e;
    LUT4 i7501_2_lut_rep_279_3_lut_4_lut (.A(\swa_swb_pwm_pulse_length_us[4] ), 
         .B(\swa_swb_pwm_pulse_length_us[3] ), .C(\swa_swb_pwm_pulse_length_us[6] ), 
         .D(\swa_swb_pwm_pulse_length_us[5] ), .Z(n52215)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;
    defparam i7501_2_lut_rep_279_3_lut_4_lut.init = 16'he000;
    LUT4 i7499_2_lut_3_lut_4_lut (.A(\swa_swb_pwm_pulse_length_us[4] ), .B(\swa_swb_pwm_pulse_length_us[3] ), 
         .C(\swa_swb_pwm_pulse_length_us[6] ), .D(\swa_swb_pwm_pulse_length_us[5] ), 
         .Z(value_out_7__N_154[6])) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B !(C)))) */ ;
    defparam i7499_2_lut_3_lut_4_lut.init = 16'h1ef0;
    LUT4 i1_2_lut (.A(\swa_swb_pwm_pulse_length_us[4] ), .B(\swa_swb_pwm_pulse_length_us[3] ), 
         .Z(value_out_7__N_154[4])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i1_2_lut.init = 16'h9999;
    LUT4 i7482_1_lut (.A(\swa_swb_pwm_pulse_length_us[3] ), .Z(value_out_7__N_154[3])) /* synthesis lut_function=(!(A)) */ ;
    defparam i7482_1_lut.init = 16'h5555;
    
endmodule
//
// Verilog Description of module pwm_reader_U2
//

module pwm_reader_U2 (state_2__N_199_c_1, us_clk, GND_net, \swa_swb_pwm_pulse_length_us[2] , 
            \swa_swb_pwm_pulse_length_us[3] , \swa_swb_pwm_pulse_length_us[4] , 
            \swa_swb_pwm_pulse_length_us[5] , \swa_swb_pwm_pulse_length_us[6] , 
            \swa_swb_pwm_pulse_length_us[7] , \swa_swb_pwm_pulse_length_us[8] , 
            \swa_swb_pwm_pulse_length_us[9] ) /* synthesis syn_module_defined=1 */ ;
    input state_2__N_199_c_1;
    input us_clk;
    input GND_net;
    output \swa_swb_pwm_pulse_length_us[2] ;
    output \swa_swb_pwm_pulse_length_us[3] ;
    output \swa_swb_pwm_pulse_length_us[4] ;
    output \swa_swb_pwm_pulse_length_us[5] ;
    output \swa_swb_pwm_pulse_length_us[6] ;
    output \swa_swb_pwm_pulse_length_us[7] ;
    output \swa_swb_pwm_pulse_length_us[8] ;
    output \swa_swb_pwm_pulse_length_us[9] ;
    
    wire us_clk /* synthesis SET_AS_NETWORK=us_clk, is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(221[10:16])
    wire [2:0]state;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(54[15:20])
    
    wire us_clk_enable_144;
    wire [15:0]time_high_count;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(57[16:31])
    
    wire n52264, n48040, n52523, n52522, n45, n12, us_clk_enable_79;
    wire [15:0]time_high_count_15__N_183;
    wire [2:0]state_2__N_180;
    
    wire n7, n51152, n52265, n4, pwm_pulse_level_flag;
    wire [15:0]time_high_count_15__N_224;
    
    wire n30718, n51050, n51051, us_clk_enable_118, n48034, n3, 
        n46781, us_clk_enable_81, n3_adj_5348, n3_adj_5349;
    wire [15:0]pwm_pulse_length_us_15__N_208;
    
    wire n9, n49002, n51156, n36411, n46641, n52373, n47135, n43901, 
        n43900, n43899, n43898, n43897, n43896, n43895, n43894, 
        n52524;
    
    LUT4 i20_4_lut_3_lut_4_lut (.A(state[1]), .B(state_2__N_199_c_1), .C(state[0]), 
         .D(state[2]), .Z(us_clk_enable_144)) /* synthesis lut_function=(A (B ((D)+!C)+!B (D))+!A !(D)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(74[13] 161[20])
    defparam i20_4_lut_3_lut_4_lut.init = 16'haa5d;
    LUT4 i1_4_lut_then_4_lut (.A(state[1]), .B(time_high_count[10]), .C(n52264), 
         .D(n48040), .Z(n52523)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_then_4_lut.init = 16'haaa8;
    LUT4 i1_4_lut_else_4_lut (.A(state[1]), .B(time_high_count[10]), .C(n52264), 
         .D(n48040), .Z(n52522)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_else_4_lut.init = 16'ha8a0;
    LUT4 i1_3_lut_4_lut (.A(time_high_count[4]), .B(n45), .C(time_high_count[3]), 
         .D(time_high_count[10]), .Z(n12)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(57[16:31])
    defparam i1_3_lut_4_lut.init = 16'h8f00;
    FD1P3AX time_high_count_i0 (.D(time_high_count_15__N_183[0]), .SP(us_clk_enable_79), 
            .CK(us_clk), .Q(time_high_count[0])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=5, LSE_RCOL=25, LSE_LLINE=159, LSE_RLINE=165 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i0.GSR = "ENABLED";
    FD1S3AX state_i0 (.D(state_2__N_180[0]), .CK(us_clk), .Q(state[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=14, LSE_LCOL=5, LSE_RCOL=25, LSE_LLINE=159, LSE_RLINE=165 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam state_i0.GSR = "ENABLED";
    LUT4 i4_4_lut_rep_328 (.A(n7), .B(time_high_count[11]), .C(time_high_count[14]), 
         .D(time_high_count[12]), .Z(n52264)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i4_4_lut_rep_328.init = 16'hfffe;
    LUT4 time_high_count_10__bdd_3_lut_40301_rep_329 (.A(time_high_count[10]), 
         .B(n51152), .C(n45), .Z(n52265)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam time_high_count_10__bdd_3_lut_40301_rep_329.init = 16'hcaca;
    LUT4 i2_4_lut (.A(state[0]), .B(state_2__N_199_c_1), .C(state[1]), 
         .D(n4), .Z(us_clk_enable_79)) /* synthesis lut_function=((B (C)+!B (C+!(D)))+!A) */ ;
    defparam i2_4_lut.init = 16'hf5f7;
    LUT4 i1_2_lut (.A(state[2]), .B(pwm_pulse_level_flag), .Z(n4)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i2_3_lut_4_lut (.A(state[1]), .B(state[2]), .C(time_high_count_15__N_224[0]), 
         .D(state[0]), .Z(time_high_count_15__N_183[0])) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i2_3_lut_4_lut.init = 16'h0020;
    LUT4 i20051_2_lut_4_lut_3_lut (.A(state[1]), .B(state[2]), .C(state[0]), 
         .Z(n30718)) /* synthesis lut_function=(A (B)+!A !(B+(C))) */ ;
    defparam i20051_2_lut_4_lut_3_lut.init = 16'h8989;
    LUT4 state_2__N_199_c_1_bdd_3_lut (.A(state_2__N_199_c_1), .B(state[1]), 
         .C(state[0]), .Z(n51050)) /* synthesis lut_function=(!(A (B)+!A (B+(C)))) */ ;
    defparam state_2__N_199_c_1_bdd_3_lut.init = 16'h2323;
    LUT4 state_2__N_199_c_1_bdd_4_lut (.A(state_2__N_199_c_1), .B(state[1]), 
         .C(state[0]), .D(pwm_pulse_level_flag), .Z(n51051)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (B+!(C (D))))) */ ;
    defparam state_2__N_199_c_1_bdd_4_lut.init = 16'h1800;
    LUT4 i39418_3_lut_rep_425 (.A(state[0]), .B(state[1]), .C(state[2]), 
         .Z(us_clk_enable_118)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;
    defparam i39418_3_lut_rep_425.init = 16'hc9c9;
    LUT4 i1_2_lut_adj_449 (.A(state[0]), .B(state[1]), .Z(n48034)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_adj_449.init = 16'h2222;
    LUT4 i1_3_lut_4_lut_adj_450 (.A(n52264), .B(time_high_count[10]), .C(time_high_count[6]), 
         .D(state[1]), .Z(n3)) /* synthesis lut_function=(A (D)+!A (B (C (D))+!B (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i1_3_lut_4_lut_adj_450.init = 16'hfb00;
    FD1S3IX state_i2 (.D(n46781), .CK(us_clk), .CD(state[2]), .Q(state[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=14, LSE_LCOL=5, LSE_RCOL=25, LSE_LLINE=159, LSE_RLINE=165 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam state_i2.GSR = "ENABLED";
    FD1S3AX state_i1 (.D(state_2__N_180[1]), .CK(us_clk), .Q(state[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=14, LSE_LCOL=5, LSE_RCOL=25, LSE_LLINE=159, LSE_RLINE=165 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam state_i1.GSR = "ENABLED";
    FD1P3AX time_high_count_i15 (.D(time_high_count_15__N_183[15]), .SP(us_clk_enable_79), 
            .CK(us_clk), .Q(time_high_count[15])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=5, LSE_RCOL=25, LSE_LLINE=159, LSE_RLINE=165 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i15.GSR = "ENABLED";
    FD1P3AX time_high_count_i14 (.D(time_high_count_15__N_183[14]), .SP(us_clk_enable_79), 
            .CK(us_clk), .Q(time_high_count[14])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=5, LSE_RCOL=25, LSE_LLINE=159, LSE_RLINE=165 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i14.GSR = "ENABLED";
    FD1P3AX time_high_count_i13 (.D(time_high_count_15__N_183[13]), .SP(us_clk_enable_79), 
            .CK(us_clk), .Q(time_high_count[13])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=5, LSE_RCOL=25, LSE_LLINE=159, LSE_RLINE=165 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i13.GSR = "ENABLED";
    FD1P3AX time_high_count_i12 (.D(time_high_count_15__N_183[12]), .SP(us_clk_enable_79), 
            .CK(us_clk), .Q(time_high_count[12])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=5, LSE_RCOL=25, LSE_LLINE=159, LSE_RLINE=165 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i12.GSR = "ENABLED";
    FD1P3AX time_high_count_i11 (.D(time_high_count_15__N_183[11]), .SP(us_clk_enable_79), 
            .CK(us_clk), .Q(time_high_count[11])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=5, LSE_RCOL=25, LSE_LLINE=159, LSE_RLINE=165 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i11.GSR = "ENABLED";
    FD1P3AX time_high_count_i10 (.D(time_high_count_15__N_183[10]), .SP(us_clk_enable_79), 
            .CK(us_clk), .Q(time_high_count[10])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=5, LSE_RCOL=25, LSE_LLINE=159, LSE_RLINE=165 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i10.GSR = "ENABLED";
    FD1P3AX time_high_count_i9 (.D(time_high_count_15__N_183[9]), .SP(us_clk_enable_79), 
            .CK(us_clk), .Q(time_high_count[9])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=5, LSE_RCOL=25, LSE_LLINE=159, LSE_RLINE=165 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i9.GSR = "ENABLED";
    FD1P3AX time_high_count_i8 (.D(time_high_count_15__N_183[8]), .SP(us_clk_enable_79), 
            .CK(us_clk), .Q(time_high_count[8])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=5, LSE_RCOL=25, LSE_LLINE=159, LSE_RLINE=165 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i8.GSR = "ENABLED";
    FD1P3AX time_high_count_i7 (.D(time_high_count_15__N_183[7]), .SP(us_clk_enable_79), 
            .CK(us_clk), .Q(time_high_count[7])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=5, LSE_RCOL=25, LSE_LLINE=159, LSE_RLINE=165 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i7.GSR = "ENABLED";
    FD1P3AX time_high_count_i6 (.D(time_high_count_15__N_183[6]), .SP(us_clk_enable_79), 
            .CK(us_clk), .Q(time_high_count[6])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=5, LSE_RCOL=25, LSE_LLINE=159, LSE_RLINE=165 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i6.GSR = "ENABLED";
    FD1P3AX time_high_count_i5 (.D(time_high_count_15__N_183[5]), .SP(us_clk_enable_79), 
            .CK(us_clk), .Q(time_high_count[5])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=5, LSE_RCOL=25, LSE_LLINE=159, LSE_RLINE=165 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i5.GSR = "ENABLED";
    FD1P3AX time_high_count_i4 (.D(time_high_count_15__N_183[4]), .SP(us_clk_enable_79), 
            .CK(us_clk), .Q(time_high_count[4])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=5, LSE_RCOL=25, LSE_LLINE=159, LSE_RLINE=165 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i4.GSR = "ENABLED";
    FD1P3AX time_high_count_i3 (.D(time_high_count_15__N_183[3]), .SP(us_clk_enable_79), 
            .CK(us_clk), .Q(time_high_count[3])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=5, LSE_RCOL=25, LSE_LLINE=159, LSE_RLINE=165 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i3.GSR = "ENABLED";
    FD1P3AX time_high_count_i2 (.D(time_high_count_15__N_183[2]), .SP(us_clk_enable_81), 
            .CK(us_clk), .Q(time_high_count[2])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=5, LSE_RCOL=25, LSE_LLINE=159, LSE_RLINE=165 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i2.GSR = "ENABLED";
    FD1P3AX time_high_count_i1 (.D(time_high_count_15__N_183[1]), .SP(us_clk_enable_81), 
            .CK(us_clk), .Q(time_high_count[1])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=5, LSE_RCOL=25, LSE_LLINE=159, LSE_RLINE=165 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i1.GSR = "ENABLED";
    LUT4 i1_3_lut_4_lut_adj_451 (.A(n52264), .B(time_high_count[10]), .C(time_high_count[7]), 
         .D(state[1]), .Z(n3_adj_5348)) /* synthesis lut_function=(A (D)+!A (B (C (D))+!B (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i1_3_lut_4_lut_adj_451.init = 16'hfb00;
    LUT4 i1_3_lut_4_lut_adj_452 (.A(n52264), .B(time_high_count[10]), .C(time_high_count[8]), 
         .D(state[1]), .Z(n3_adj_5349)) /* synthesis lut_function=(A (D)+!A (B (C (D))+!B (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i1_3_lut_4_lut_adj_452.init = 16'hfb00;
    LUT4 i1_2_lut_3_lut (.A(n52264), .B(time_high_count[10]), .C(time_high_count[9]), 
         .Z(pwm_pulse_length_us_15__N_208[9])) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i1_2_lut_3_lut.init = 16'hfbfb;
    LUT4 n45_bdd_4_lut_40300 (.A(time_high_count[10]), .B(time_high_count[4]), 
         .C(time_high_count[5]), .D(time_high_count[3]), .Z(n51152)) /* synthesis lut_function=(!(A (B+(C))+!A !(B (C)+!B (C (D))))) */ ;
    defparam n45_bdd_4_lut_40300.init = 16'h5242;
    LUT4 i3_4_lut (.A(time_high_count[6]), .B(time_high_count[8]), .C(time_high_count[9]), 
         .D(time_high_count[7]), .Z(n45)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(57[16:31])
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i2_2_lut (.A(time_high_count[13]), .B(time_high_count[15]), .Z(n7)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i3_4_lut_4_lut (.A(n52264), .B(n12), .C(n9), .D(state[1]), 
         .Z(n49002)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i3_4_lut_4_lut.init = 16'h0100;
    LUT4 gnd_bdd_2_lut_40274_3_lut_4_lut (.A(n52265), .B(state[1]), .C(time_high_count[2]), 
         .D(n52264), .Z(n51156)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam gnd_bdd_2_lut_40274_3_lut_4_lut.init = 16'h0080;
    LUT4 i1_4_lut (.A(time_high_count[4]), .B(n48040), .C(time_high_count[10]), 
         .D(time_high_count[3]), .Z(n9)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(57[16:31])
    defparam i1_4_lut.init = 16'hc0c8;
    LUT4 i1_2_lut_adj_453 (.A(n45), .B(time_high_count[5]), .Z(n48040)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_453.init = 16'h8888;
    LUT4 i39617_4_lut (.A(n52264), .B(time_high_count[5]), .C(time_high_count[10]), 
         .D(n45), .Z(pwm_pulse_length_us_15__N_208[5])) /* synthesis lut_function=(!(A+(B (C (D))+!B (C)))) */ ;
    defparam i39617_4_lut.init = 16'h0545;
    LUT4 i1_2_lut_4_lut_4_lut (.A(state[0]), .B(time_high_count_15__N_224[9]), 
         .C(state[1]), .D(state[2]), .Z(time_high_count_15__N_183[9])) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut.init = 16'h0040;
    LUT4 i1_2_lut_4_lut_4_lut_adj_454 (.A(state[0]), .B(time_high_count_15__N_224[15]), 
         .C(state[1]), .D(state[2]), .Z(time_high_count_15__N_183[15])) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_454.init = 16'h0040;
    LUT4 i1_2_lut_4_lut_4_lut_adj_455 (.A(state[0]), .B(time_high_count_15__N_224[11]), 
         .C(state[1]), .D(state[2]), .Z(time_high_count_15__N_183[11])) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_455.init = 16'h0040;
    LUT4 i1_2_lut_4_lut_4_lut_adj_456 (.A(state[0]), .B(time_high_count_15__N_224[1]), 
         .C(state[1]), .D(state[2]), .Z(time_high_count_15__N_183[1])) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_456.init = 16'h0040;
    LUT4 i1_2_lut_4_lut_4_lut_adj_457 (.A(state[0]), .B(time_high_count_15__N_224[2]), 
         .C(state[1]), .D(state[2]), .Z(time_high_count_15__N_183[2])) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_457.init = 16'h0040;
    LUT4 i1_2_lut_4_lut_4_lut_adj_458 (.A(state[0]), .B(time_high_count_15__N_224[10]), 
         .C(state[1]), .D(state[2]), .Z(time_high_count_15__N_183[10])) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_458.init = 16'h0040;
    PFUMX i40203 (.BLUT(n51051), .ALUT(n51050), .C0(state[2]), .Z(state_2__N_180[1]));
    LUT4 i1_2_lut_4_lut_4_lut_adj_459 (.A(state[0]), .B(time_high_count_15__N_224[3]), 
         .C(state[1]), .D(state[2]), .Z(time_high_count_15__N_183[3])) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_459.init = 16'h0040;
    LUT4 i1_2_lut_4_lut_4_lut_adj_460 (.A(state[0]), .B(time_high_count_15__N_224[4]), 
         .C(state[1]), .D(state[2]), .Z(time_high_count_15__N_183[4])) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_460.init = 16'h0040;
    LUT4 i1_2_lut_4_lut_4_lut_adj_461 (.A(state[0]), .B(time_high_count_15__N_224[14]), 
         .C(state[1]), .D(state[2]), .Z(time_high_count_15__N_183[14])) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_461.init = 16'h0040;
    LUT4 i1_2_lut_4_lut_4_lut_adj_462 (.A(state[0]), .B(time_high_count_15__N_224[5]), 
         .C(state[1]), .D(state[2]), .Z(time_high_count_15__N_183[5])) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_462.init = 16'h0040;
    LUT4 i1_2_lut_4_lut_4_lut_adj_463 (.A(state[0]), .B(time_high_count_15__N_224[13]), 
         .C(state[1]), .D(state[2]), .Z(time_high_count_15__N_183[13])) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_463.init = 16'h0040;
    LUT4 i1_2_lut_4_lut_4_lut_adj_464 (.A(state[0]), .B(time_high_count_15__N_224[8]), 
         .C(state[1]), .D(state[2]), .Z(time_high_count_15__N_183[8])) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_464.init = 16'h0040;
    LUT4 i1_2_lut_4_lut_4_lut_adj_465 (.A(state[0]), .B(time_high_count_15__N_224[6]), 
         .C(state[1]), .D(state[2]), .Z(time_high_count_15__N_183[6])) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_465.init = 16'h0040;
    LUT4 i1_2_lut_4_lut_4_lut_adj_466 (.A(state[0]), .B(time_high_count_15__N_224[7]), 
         .C(state[1]), .D(state[2]), .Z(time_high_count_15__N_183[7])) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_466.init = 16'h0040;
    LUT4 i1_2_lut_4_lut_4_lut_adj_467 (.A(state[0]), .B(time_high_count_15__N_224[12]), 
         .C(state[1]), .D(state[2]), .Z(time_high_count_15__N_183[12])) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i1_2_lut_4_lut_4_lut_adj_467.init = 16'h0040;
    LUT4 i25790_2_lut (.A(state[2]), .B(state[1]), .Z(n36411)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i25790_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_468 (.A(pwm_pulse_level_flag), .B(state[1]), .C(state_2__N_199_c_1), 
         .D(state[0]), .Z(n46641)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(74[13] 161[20])
    defparam i1_4_lut_adj_468.init = 16'heccc;
    LUT4 state_2__N_199_c_1_bdd_4_lut_40202 (.A(state_2__N_199_c_1), .B(state[2]), 
         .C(state[0]), .D(state[1]), .Z(state_2__N_180[0])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B ((D)+!C)))) */ ;
    defparam state_2__N_199_c_1_bdd_4_lut_40202.init = 16'h3173;
    LUT4 i21_4_lut (.A(state_2__N_199_c_1), .B(pwm_pulse_level_flag), .C(state[1]), 
         .D(state[0]), .Z(n46781)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A ((D)+!C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(74[13] 161[20])
    defparam i21_4_lut.init = 16'h0a70;
    LUT4 i39935_4_lut (.A(pwm_pulse_level_flag), .B(n48034), .C(state_2__N_199_c_1), 
         .D(state[2]), .Z(us_clk_enable_81)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))))) */ ;
    defparam i39935_4_lut.init = 16'h3337;
    LUT4 pwm_pulse_level_flag_I_0_55_1_lut_rep_437 (.A(pwm_pulse_level_flag), 
         .Z(n52373)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[46:74])
    defparam pwm_pulse_level_flag_I_0_55_1_lut_rep_437.init = 16'h5555;
    LUT4 i1_2_lut_2_lut (.A(pwm_pulse_level_flag), .B(state_2__N_199_c_1), 
         .Z(n47135)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[46:74])
    defparam i1_2_lut_2_lut.init = 16'h4444;
    CCU2D add_3759_17 (.A0(n52373), .B0(state_2__N_199_c_1), .C0(time_high_count[15]), 
          .D0(pwm_pulse_level_flag), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43901), .S0(time_high_count_15__N_224[15]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3759_17.INIT0 = 16'hf070;
    defparam add_3759_17.INIT1 = 16'h0000;
    defparam add_3759_17.INJECT1_0 = "NO";
    defparam add_3759_17.INJECT1_1 = "NO";
    CCU2D add_3759_15 (.A0(n52373), .B0(state_2__N_199_c_1), .C0(time_high_count[13]), 
          .D0(pwm_pulse_level_flag), .A1(n52373), .B1(state_2__N_199_c_1), 
          .C1(time_high_count[14]), .D1(pwm_pulse_level_flag), .CIN(n43900), 
          .COUT(n43901), .S0(time_high_count_15__N_224[13]), .S1(time_high_count_15__N_224[14]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3759_15.INIT0 = 16'hf070;
    defparam add_3759_15.INIT1 = 16'hf070;
    defparam add_3759_15.INJECT1_0 = "NO";
    defparam add_3759_15.INJECT1_1 = "NO";
    CCU2D add_3759_13 (.A0(n52373), .B0(state_2__N_199_c_1), .C0(time_high_count[11]), 
          .D0(pwm_pulse_level_flag), .A1(n52373), .B1(state_2__N_199_c_1), 
          .C1(time_high_count[12]), .D1(pwm_pulse_level_flag), .CIN(n43899), 
          .COUT(n43900), .S0(time_high_count_15__N_224[11]), .S1(time_high_count_15__N_224[12]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3759_13.INIT0 = 16'hf070;
    defparam add_3759_13.INIT1 = 16'hf070;
    defparam add_3759_13.INJECT1_0 = "NO";
    defparam add_3759_13.INJECT1_1 = "NO";
    CCU2D add_3759_11 (.A0(n52373), .B0(state_2__N_199_c_1), .C0(time_high_count[9]), 
          .D0(pwm_pulse_level_flag), .A1(n52373), .B1(state_2__N_199_c_1), 
          .C1(time_high_count[10]), .D1(pwm_pulse_level_flag), .CIN(n43898), 
          .COUT(n43899), .S0(time_high_count_15__N_224[9]), .S1(time_high_count_15__N_224[10]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3759_11.INIT0 = 16'hf070;
    defparam add_3759_11.INIT1 = 16'hf070;
    defparam add_3759_11.INJECT1_0 = "NO";
    defparam add_3759_11.INJECT1_1 = "NO";
    CCU2D add_3759_9 (.A0(n52373), .B0(state_2__N_199_c_1), .C0(time_high_count[7]), 
          .D0(pwm_pulse_level_flag), .A1(n52373), .B1(state_2__N_199_c_1), 
          .C1(time_high_count[8]), .D1(pwm_pulse_level_flag), .CIN(n43897), 
          .COUT(n43898), .S0(time_high_count_15__N_224[7]), .S1(time_high_count_15__N_224[8]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3759_9.INIT0 = 16'hf070;
    defparam add_3759_9.INIT1 = 16'hf070;
    defparam add_3759_9.INJECT1_0 = "NO";
    defparam add_3759_9.INJECT1_1 = "NO";
    CCU2D add_3759_7 (.A0(n52373), .B0(state_2__N_199_c_1), .C0(time_high_count[5]), 
          .D0(pwm_pulse_level_flag), .A1(n52373), .B1(state_2__N_199_c_1), 
          .C1(time_high_count[6]), .D1(pwm_pulse_level_flag), .CIN(n43896), 
          .COUT(n43897), .S0(time_high_count_15__N_224[5]), .S1(time_high_count_15__N_224[6]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3759_7.INIT0 = 16'hf070;
    defparam add_3759_7.INIT1 = 16'hf070;
    defparam add_3759_7.INJECT1_0 = "NO";
    defparam add_3759_7.INJECT1_1 = "NO";
    CCU2D add_3759_5 (.A0(n52373), .B0(state_2__N_199_c_1), .C0(time_high_count[3]), 
          .D0(pwm_pulse_level_flag), .A1(n52373), .B1(state_2__N_199_c_1), 
          .C1(time_high_count[4]), .D1(pwm_pulse_level_flag), .CIN(n43895), 
          .COUT(n43896), .S0(time_high_count_15__N_224[3]), .S1(time_high_count_15__N_224[4]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3759_5.INIT0 = 16'hf070;
    defparam add_3759_5.INIT1 = 16'hf070;
    defparam add_3759_5.INJECT1_0 = "NO";
    defparam add_3759_5.INJECT1_1 = "NO";
    CCU2D add_3759_3 (.A0(n52373), .B0(state_2__N_199_c_1), .C0(time_high_count[1]), 
          .D0(pwm_pulse_level_flag), .A1(n52373), .B1(state_2__N_199_c_1), 
          .C1(time_high_count[2]), .D1(pwm_pulse_level_flag), .CIN(n43894), 
          .COUT(n43895), .S0(time_high_count_15__N_224[1]), .S1(time_high_count_15__N_224[2]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3759_3.INIT0 = 16'hf070;
    defparam add_3759_3.INIT1 = 16'hf070;
    defparam add_3759_3.INJECT1_0 = "NO";
    defparam add_3759_3.INJECT1_1 = "NO";
    CCU2D add_3759_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(time_high_count[0]), .B1(n47135), .C1(state_2__N_199_c_1), 
          .D1(pwm_pulse_level_flag), .COUT(n43894), .S1(time_high_count_15__N_224[0]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3759_1.INIT0 = 16'hF000;
    defparam add_3759_1.INIT1 = 16'hd222;
    defparam add_3759_1.INJECT1_0 = "NO";
    defparam add_3759_1.INJECT1_1 = "NO";
    PFUMX i40942 (.BLUT(n52522), .ALUT(n52523), .C0(time_high_count[4]), 
          .Z(n52524));
    FD1P3JX time_high_us_i2 (.D(n51156), .SP(us_clk_enable_118), .PD(n30718), 
            .CK(us_clk), .Q(\swa_swb_pwm_pulse_length_us[2] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=5, LSE_RCOL=25, LSE_LLINE=159, LSE_RLINE=165 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i2.GSR = "ENABLED";
    FD1P3JX time_high_us_i3 (.D(n49002), .SP(us_clk_enable_118), .PD(n30718), 
            .CK(us_clk), .Q(\swa_swb_pwm_pulse_length_us[3] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=5, LSE_RCOL=25, LSE_LLINE=159, LSE_RLINE=165 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i3.GSR = "ENABLED";
    FD1P3JX time_high_us_i4 (.D(n52524), .SP(us_clk_enable_118), .PD(n30718), 
            .CK(us_clk), .Q(\swa_swb_pwm_pulse_length_us[4] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=5, LSE_RCOL=25, LSE_LLINE=159, LSE_RLINE=165 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i4.GSR = "ENABLED";
    FD1P3IX time_high_us_i5 (.D(pwm_pulse_length_us_15__N_208[5]), .SP(us_clk_enable_118), 
            .CD(n30718), .CK(us_clk), .Q(\swa_swb_pwm_pulse_length_us[5] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=5, LSE_RCOL=25, LSE_LLINE=159, LSE_RLINE=165 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i5.GSR = "ENABLED";
    FD1P3JX time_high_us_i6 (.D(n3), .SP(us_clk_enable_118), .PD(n30718), 
            .CK(us_clk), .Q(\swa_swb_pwm_pulse_length_us[6] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=5, LSE_RCOL=25, LSE_LLINE=159, LSE_RLINE=165 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i6.GSR = "ENABLED";
    FD1P3JX time_high_us_i7 (.D(n3_adj_5348), .SP(us_clk_enable_118), .PD(n30718), 
            .CK(us_clk), .Q(\swa_swb_pwm_pulse_length_us[7] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=5, LSE_RCOL=25, LSE_LLINE=159, LSE_RLINE=165 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i7.GSR = "ENABLED";
    FD1P3JX time_high_us_i8 (.D(n3_adj_5349), .SP(us_clk_enable_118), .PD(n30718), 
            .CK(us_clk), .Q(\swa_swb_pwm_pulse_length_us[8] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=5, LSE_RCOL=25, LSE_LLINE=159, LSE_RLINE=165 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i8.GSR = "ENABLED";
    FD1P3IX time_high_us_i9 (.D(pwm_pulse_length_us_15__N_208[9]), .SP(us_clk_enable_118), 
            .CD(n30718), .CK(us_clk), .Q(\swa_swb_pwm_pulse_length_us[9] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=5, LSE_RCOL=25, LSE_LLINE=159, LSE_RLINE=165 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i9.GSR = "ENABLED";
    FD1P3IX pwm_pulse_level_flag_46 (.D(n46641), .SP(us_clk_enable_144), 
            .CD(n36411), .CK(us_clk), .Q(pwm_pulse_level_flag)) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=5, LSE_RCOL=25, LSE_LLINE=159, LSE_RLINE=165 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam pwm_pulse_level_flag_46.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module pwm_reader_U3
//

module pwm_reader_U3 (state_2__N_199_c_1, us_clk, GND_net, \roll_pwm_pulse_length_us[2] , 
            \roll_pwm_pulse_length_us[3] , \roll_pwm_pulse_length_us[4] , 
            \roll_pwm_pulse_length_us[5] , \roll_pwm_pulse_length_us[6] , 
            \roll_pwm_pulse_length_us[7] , \roll_pwm_pulse_length_us[8] , 
            \roll_pwm_pulse_length_us[9] ) /* synthesis syn_module_defined=1 */ ;
    input state_2__N_199_c_1;
    input us_clk;
    input GND_net;
    output \roll_pwm_pulse_length_us[2] ;
    output \roll_pwm_pulse_length_us[3] ;
    output \roll_pwm_pulse_length_us[4] ;
    output \roll_pwm_pulse_length_us[5] ;
    output \roll_pwm_pulse_length_us[6] ;
    output \roll_pwm_pulse_length_us[7] ;
    output \roll_pwm_pulse_length_us[8] ;
    output \roll_pwm_pulse_length_us[9] ;
    
    wire us_clk /* synthesis SET_AS_NETWORK=us_clk, is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(221[10:16])
    wire [2:0]state;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(54[15:20])
    
    wire us_clk_enable_146;
    wire [15:0]time_high_count;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(57[16:31])
    
    wire n35428, n48043, n52516, n45, n12, us_clk_enable_38;
    wire [15:0]time_high_count_15__N_183;
    wire [2:0]state_2__N_180;
    
    wire n51094, n52278, n4, pwm_pulse_level_flag, n46787, us_clk_enable_40, 
        n51031, n51032, n3, n3_adj_5346, n3_adj_5347, n52392, n47131;
    wire [15:0]pwm_pulse_length_us_15__N_208;
    
    wire n47951, n52517, n7, n9, n48998, us_clk_enable_134, n51098, 
        n36401, n46549;
    wire [15:0]time_high_count_15__N_224;
    
    wire n30680, n43933, n43932, n43931, n43930, n43929, n43928, 
        n43927, n43926, n52518;
    
    LUT4 i20_4_lut_3_lut_4_lut (.A(state[1]), .B(state_2__N_199_c_1), .C(state[0]), 
         .D(state[2]), .Z(us_clk_enable_146)) /* synthesis lut_function=(A (B ((D)+!C)+!B (D))+!A !(D)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i20_4_lut_3_lut_4_lut.init = 16'haa5d;
    LUT4 i1_4_lut_else_4_lut (.A(state[1]), .B(time_high_count[10]), .C(n35428), 
         .D(n48043), .Z(n52516)) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;
    defparam i1_4_lut_else_4_lut.init = 16'ha8a0;
    LUT4 i1_3_lut_4_lut (.A(time_high_count[4]), .B(n45), .C(time_high_count[3]), 
         .D(time_high_count[10]), .Z(n12)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(57[16:31])
    defparam i1_3_lut_4_lut.init = 16'h8f00;
    FD1P3AX time_high_count_i0 (.D(time_high_count_15__N_183[0]), .SP(us_clk_enable_38), 
            .CK(us_clk), .Q(time_high_count[0])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=52, LSE_RCOL=25, LSE_LLINE=92, LSE_RLINE=98 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i0.GSR = "ENABLED";
    FD1S3AX state_i0 (.D(state_2__N_180[0]), .CK(us_clk), .Q(state[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=14, LSE_LCOL=52, LSE_RCOL=25, LSE_LLINE=92, LSE_RLINE=98 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam state_i0.GSR = "ENABLED";
    LUT4 time_high_count_10__bdd_3_lut_40426_rep_342 (.A(time_high_count[10]), 
         .B(n51094), .C(n45), .Z(n52278)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam time_high_count_10__bdd_3_lut_40426_rep_342.init = 16'hcaca;
    LUT4 i2_4_lut (.A(state[0]), .B(state_2__N_199_c_1), .C(state[1]), 
         .D(n4), .Z(us_clk_enable_38)) /* synthesis lut_function=((B (C)+!B (C+!(D)))+!A) */ ;
    defparam i2_4_lut.init = 16'hf5f7;
    LUT4 i1_2_lut (.A(state[2]), .B(pwm_pulse_level_flag), .Z(n4)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    FD1S3IX state_i2 (.D(n46787), .CK(us_clk), .CD(state[2]), .Q(state[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=14, LSE_LCOL=52, LSE_RCOL=25, LSE_LLINE=92, LSE_RLINE=98 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam state_i2.GSR = "ENABLED";
    FD1S3AX state_i1 (.D(state_2__N_180[1]), .CK(us_clk), .Q(state[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=14, LSE_LCOL=52, LSE_RCOL=25, LSE_LLINE=92, LSE_RLINE=98 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam state_i1.GSR = "ENABLED";
    FD1P3AX time_high_count_i15 (.D(time_high_count_15__N_183[15]), .SP(us_clk_enable_38), 
            .CK(us_clk), .Q(time_high_count[15])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=52, LSE_RCOL=25, LSE_LLINE=92, LSE_RLINE=98 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i15.GSR = "ENABLED";
    FD1P3AX time_high_count_i14 (.D(time_high_count_15__N_183[14]), .SP(us_clk_enable_38), 
            .CK(us_clk), .Q(time_high_count[14])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=52, LSE_RCOL=25, LSE_LLINE=92, LSE_RLINE=98 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i14.GSR = "ENABLED";
    FD1P3AX time_high_count_i13 (.D(time_high_count_15__N_183[13]), .SP(us_clk_enable_38), 
            .CK(us_clk), .Q(time_high_count[13])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=52, LSE_RCOL=25, LSE_LLINE=92, LSE_RLINE=98 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i13.GSR = "ENABLED";
    FD1P3AX time_high_count_i12 (.D(time_high_count_15__N_183[12]), .SP(us_clk_enable_38), 
            .CK(us_clk), .Q(time_high_count[12])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=52, LSE_RCOL=25, LSE_LLINE=92, LSE_RLINE=98 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i12.GSR = "ENABLED";
    FD1P3AX time_high_count_i11 (.D(time_high_count_15__N_183[11]), .SP(us_clk_enable_38), 
            .CK(us_clk), .Q(time_high_count[11])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=52, LSE_RCOL=25, LSE_LLINE=92, LSE_RLINE=98 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i11.GSR = "ENABLED";
    FD1P3AX time_high_count_i10 (.D(time_high_count_15__N_183[10]), .SP(us_clk_enable_38), 
            .CK(us_clk), .Q(time_high_count[10])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=52, LSE_RCOL=25, LSE_LLINE=92, LSE_RLINE=98 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i10.GSR = "ENABLED";
    FD1P3AX time_high_count_i9 (.D(time_high_count_15__N_183[9]), .SP(us_clk_enable_38), 
            .CK(us_clk), .Q(time_high_count[9])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=52, LSE_RCOL=25, LSE_LLINE=92, LSE_RLINE=98 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i9.GSR = "ENABLED";
    FD1P3AX time_high_count_i8 (.D(time_high_count_15__N_183[8]), .SP(us_clk_enable_38), 
            .CK(us_clk), .Q(time_high_count[8])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=52, LSE_RCOL=25, LSE_LLINE=92, LSE_RLINE=98 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i8.GSR = "ENABLED";
    FD1P3AX time_high_count_i7 (.D(time_high_count_15__N_183[7]), .SP(us_clk_enable_38), 
            .CK(us_clk), .Q(time_high_count[7])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=52, LSE_RCOL=25, LSE_LLINE=92, LSE_RLINE=98 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i7.GSR = "ENABLED";
    FD1P3AX time_high_count_i6 (.D(time_high_count_15__N_183[6]), .SP(us_clk_enable_38), 
            .CK(us_clk), .Q(time_high_count[6])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=52, LSE_RCOL=25, LSE_LLINE=92, LSE_RLINE=98 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i6.GSR = "ENABLED";
    FD1P3AX time_high_count_i5 (.D(time_high_count_15__N_183[5]), .SP(us_clk_enable_38), 
            .CK(us_clk), .Q(time_high_count[5])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=52, LSE_RCOL=25, LSE_LLINE=92, LSE_RLINE=98 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i5.GSR = "ENABLED";
    FD1P3AX time_high_count_i4 (.D(time_high_count_15__N_183[4]), .SP(us_clk_enable_38), 
            .CK(us_clk), .Q(time_high_count[4])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=52, LSE_RCOL=25, LSE_LLINE=92, LSE_RLINE=98 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i4.GSR = "ENABLED";
    FD1P3AX time_high_count_i3 (.D(time_high_count_15__N_183[3]), .SP(us_clk_enable_38), 
            .CK(us_clk), .Q(time_high_count[3])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=52, LSE_RCOL=25, LSE_LLINE=92, LSE_RLINE=98 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i3.GSR = "ENABLED";
    FD1P3AX time_high_count_i2 (.D(time_high_count_15__N_183[2]), .SP(us_clk_enable_40), 
            .CK(us_clk), .Q(time_high_count[2])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=52, LSE_RCOL=25, LSE_LLINE=92, LSE_RLINE=98 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i2.GSR = "ENABLED";
    FD1P3AX time_high_count_i1 (.D(time_high_count_15__N_183[1]), .SP(us_clk_enable_40), 
            .CK(us_clk), .Q(time_high_count[1])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=52, LSE_RCOL=25, LSE_LLINE=92, LSE_RLINE=98 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i1.GSR = "ENABLED";
    LUT4 state_1__bdd_3_lut (.A(state[1]), .B(state[0]), .C(state_2__N_199_c_1), 
         .Z(n51031)) /* synthesis lut_function=(!(A+!((C)+!B))) */ ;
    defparam state_1__bdd_3_lut.init = 16'h5151;
    LUT4 state_1__bdd_4_lut_40219 (.A(state[1]), .B(pwm_pulse_level_flag), 
         .C(state[0]), .D(state_2__N_199_c_1), .Z(n51032)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (((D)+!C)+!B))) */ ;
    defparam state_1__bdd_4_lut_40219.init = 16'h0840;
    LUT4 state_0__bdd_4_lut (.A(state[0]), .B(state[2]), .C(state[1]), 
         .D(state_2__N_199_c_1), .Z(state_2__N_180[0])) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B+(C (D))))) */ ;
    defparam state_0__bdd_4_lut.init = 16'h233b;
    LUT4 i1_3_lut_4_lut_adj_428 (.A(n35428), .B(time_high_count[10]), .C(time_high_count[6]), 
         .D(state[1]), .Z(n3)) /* synthesis lut_function=(A (D)+!A (B (C (D))+!B (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i1_3_lut_4_lut_adj_428.init = 16'hfb00;
    LUT4 i1_3_lut_4_lut_adj_429 (.A(n35428), .B(time_high_count[10]), .C(time_high_count[7]), 
         .D(state[1]), .Z(n3_adj_5346)) /* synthesis lut_function=(A (D)+!A (B (C (D))+!B (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i1_3_lut_4_lut_adj_429.init = 16'hfb00;
    LUT4 i1_3_lut_4_lut_adj_430 (.A(n35428), .B(time_high_count[10]), .C(time_high_count[8]), 
         .D(state[1]), .Z(n3_adj_5347)) /* synthesis lut_function=(A (D)+!A (B (C (D))+!B (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i1_3_lut_4_lut_adj_430.init = 16'hfb00;
    LUT4 n45_bdd_4_lut_40425 (.A(time_high_count[10]), .B(time_high_count[4]), 
         .C(time_high_count[5]), .D(time_high_count[3]), .Z(n51094)) /* synthesis lut_function=(!(A (B+(C))+!A !(B (C)+!B (C (D))))) */ ;
    defparam n45_bdd_4_lut_40425.init = 16'h5242;
    LUT4 pwm_pulse_level_flag_I_0_55_1_lut_rep_456 (.A(pwm_pulse_level_flag), 
         .Z(n52392)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[46:74])
    defparam pwm_pulse_level_flag_I_0_55_1_lut_rep_456.init = 16'h5555;
    LUT4 i1_2_lut_2_lut (.A(pwm_pulse_level_flag), .B(state_2__N_199_c_1), 
         .Z(n47131)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[46:74])
    defparam i1_2_lut_2_lut.init = 16'h4444;
    LUT4 i1_2_lut_3_lut (.A(n35428), .B(time_high_count[10]), .C(time_high_count[9]), 
         .Z(pwm_pulse_length_us_15__N_208[9])) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i1_2_lut_3_lut.init = 16'hfbfb;
    LUT4 i21_4_lut (.A(state_2__N_199_c_1), .B(pwm_pulse_level_flag), .C(state[1]), 
         .D(state[0]), .Z(n46787)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A ((D)+!C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(74[13] 161[20])
    defparam i21_4_lut.init = 16'h0a70;
    LUT4 i39709_4_lut (.A(pwm_pulse_level_flag), .B(n47951), .C(state_2__N_199_c_1), 
         .D(state[2]), .Z(us_clk_enable_40)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))))) */ ;
    defparam i39709_4_lut.init = 16'h3337;
    LUT4 i1_2_lut_adj_431 (.A(state[0]), .B(state[1]), .Z(n47951)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i1_2_lut_adj_431.init = 16'h2222;
    LUT4 i1_4_lut_then_4_lut (.A(state[1]), .B(time_high_count[10]), .C(n35428), 
         .D(n48043), .Z(n52517)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i1_4_lut_then_4_lut.init = 16'haaa8;
    LUT4 i4_4_lut (.A(n7), .B(time_high_count[14]), .C(time_high_count[12]), 
         .D(time_high_count[11]), .Z(n35428)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i4_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut (.A(time_high_count[15]), .B(time_high_count[13]), .Z(n7)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i3_4_lut (.A(time_high_count[9]), .B(time_high_count[8]), .C(time_high_count[7]), 
         .D(time_high_count[6]), .Z(n45)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(57[16:31])
    defparam i3_4_lut.init = 16'h8000;
    LUT4 i3_4_lut_adj_432 (.A(state[1]), .B(n9), .C(n35428), .D(n12), 
         .Z(n48998)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i3_4_lut_adj_432.init = 16'h0002;
    LUT4 i1_4_lut (.A(time_high_count[4]), .B(n48043), .C(time_high_count[10]), 
         .D(time_high_count[3]), .Z(n9)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(57[16:31])
    defparam i1_4_lut.init = 16'hc0c8;
    LUT4 i1_2_lut_adj_433 (.A(n45), .B(time_high_count[5]), .Z(n48043)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_adj_433.init = 16'h8888;
    LUT4 i39607_4_lut (.A(n35428), .B(time_high_count[5]), .C(time_high_count[10]), 
         .D(n45), .Z(pwm_pulse_length_us_15__N_208[5])) /* synthesis lut_function=(!(A+(B (C (D))+!B (C)))) */ ;
    defparam i39607_4_lut.init = 16'h0545;
    LUT4 i39416_3_lut_rep_417 (.A(state[0]), .B(state[1]), .C(state[2]), 
         .Z(us_clk_enable_134)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;
    defparam i39416_3_lut_rep_417.init = 16'hc9c9;
    LUT4 gnd_bdd_2_lut_40228_3_lut_4_lut (.A(n52278), .B(state[1]), .C(time_high_count[2]), 
         .D(n35428), .Z(n51098)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam gnd_bdd_2_lut_40228_3_lut_4_lut.init = 16'h0080;
    PFUMX i40188 (.BLUT(n51032), .ALUT(n51031), .C0(state[2]), .Z(state_2__N_180[1]));
    LUT4 i25780_2_lut (.A(state[2]), .B(state[1]), .Z(n36401)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i25780_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_434 (.A(pwm_pulse_level_flag), .B(state[1]), .C(state_2__N_199_c_1), 
         .D(state[0]), .Z(n46549)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(74[13] 161[20])
    defparam i1_4_lut_adj_434.init = 16'heccc;
    LUT4 i2_3_lut_4_lut (.A(state[1]), .B(state[2]), .C(time_high_count_15__N_224[0]), 
         .D(state[0]), .Z(time_high_count_15__N_183[0])) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i2_3_lut_4_lut.init = 16'h0020;
    LUT4 i20013_2_lut_4_lut_3_lut (.A(state[1]), .B(state[2]), .C(state[0]), 
         .Z(n30680)) /* synthesis lut_function=(A (B)+!A !(B+(C))) */ ;
    defparam i20013_2_lut_4_lut_3_lut.init = 16'h8989;
    CCU2D add_3751_17 (.A0(n52392), .B0(state_2__N_199_c_1), .C0(time_high_count[15]), 
          .D0(pwm_pulse_level_flag), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43933), .S0(time_high_count_15__N_224[15]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3751_17.INIT0 = 16'hf070;
    defparam add_3751_17.INIT1 = 16'h0000;
    defparam add_3751_17.INJECT1_0 = "NO";
    defparam add_3751_17.INJECT1_1 = "NO";
    CCU2D add_3751_15 (.A0(n52392), .B0(state_2__N_199_c_1), .C0(time_high_count[13]), 
          .D0(pwm_pulse_level_flag), .A1(n52392), .B1(state_2__N_199_c_1), 
          .C1(time_high_count[14]), .D1(pwm_pulse_level_flag), .CIN(n43932), 
          .COUT(n43933), .S0(time_high_count_15__N_224[13]), .S1(time_high_count_15__N_224[14]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3751_15.INIT0 = 16'hf070;
    defparam add_3751_15.INIT1 = 16'hf070;
    defparam add_3751_15.INJECT1_0 = "NO";
    defparam add_3751_15.INJECT1_1 = "NO";
    CCU2D add_3751_13 (.A0(n52392), .B0(state_2__N_199_c_1), .C0(time_high_count[11]), 
          .D0(pwm_pulse_level_flag), .A1(n52392), .B1(state_2__N_199_c_1), 
          .C1(time_high_count[12]), .D1(pwm_pulse_level_flag), .CIN(n43931), 
          .COUT(n43932), .S0(time_high_count_15__N_224[11]), .S1(time_high_count_15__N_224[12]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3751_13.INIT0 = 16'hf070;
    defparam add_3751_13.INIT1 = 16'hf070;
    defparam add_3751_13.INJECT1_0 = "NO";
    defparam add_3751_13.INJECT1_1 = "NO";
    CCU2D add_3751_11 (.A0(n52392), .B0(state_2__N_199_c_1), .C0(time_high_count[9]), 
          .D0(pwm_pulse_level_flag), .A1(n52392), .B1(state_2__N_199_c_1), 
          .C1(time_high_count[10]), .D1(pwm_pulse_level_flag), .CIN(n43930), 
          .COUT(n43931), .S0(time_high_count_15__N_224[9]), .S1(time_high_count_15__N_224[10]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3751_11.INIT0 = 16'hf070;
    defparam add_3751_11.INIT1 = 16'hf070;
    defparam add_3751_11.INJECT1_0 = "NO";
    defparam add_3751_11.INJECT1_1 = "NO";
    CCU2D add_3751_9 (.A0(n52392), .B0(state_2__N_199_c_1), .C0(time_high_count[7]), 
          .D0(pwm_pulse_level_flag), .A1(n52392), .B1(state_2__N_199_c_1), 
          .C1(time_high_count[8]), .D1(pwm_pulse_level_flag), .CIN(n43929), 
          .COUT(n43930), .S0(time_high_count_15__N_224[7]), .S1(time_high_count_15__N_224[8]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3751_9.INIT0 = 16'hf070;
    defparam add_3751_9.INIT1 = 16'hf070;
    defparam add_3751_9.INJECT1_0 = "NO";
    defparam add_3751_9.INJECT1_1 = "NO";
    CCU2D add_3751_7 (.A0(n52392), .B0(state_2__N_199_c_1), .C0(time_high_count[5]), 
          .D0(pwm_pulse_level_flag), .A1(n52392), .B1(state_2__N_199_c_1), 
          .C1(time_high_count[6]), .D1(pwm_pulse_level_flag), .CIN(n43928), 
          .COUT(n43929), .S0(time_high_count_15__N_224[5]), .S1(time_high_count_15__N_224[6]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3751_7.INIT0 = 16'hf070;
    defparam add_3751_7.INIT1 = 16'hf070;
    defparam add_3751_7.INJECT1_0 = "NO";
    defparam add_3751_7.INJECT1_1 = "NO";
    CCU2D add_3751_5 (.A0(n52392), .B0(state_2__N_199_c_1), .C0(time_high_count[3]), 
          .D0(pwm_pulse_level_flag), .A1(n52392), .B1(state_2__N_199_c_1), 
          .C1(time_high_count[4]), .D1(pwm_pulse_level_flag), .CIN(n43927), 
          .COUT(n43928), .S0(time_high_count_15__N_224[3]), .S1(time_high_count_15__N_224[4]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3751_5.INIT0 = 16'hf070;
    defparam add_3751_5.INIT1 = 16'hf070;
    defparam add_3751_5.INJECT1_0 = "NO";
    defparam add_3751_5.INJECT1_1 = "NO";
    CCU2D add_3751_3 (.A0(n52392), .B0(state_2__N_199_c_1), .C0(time_high_count[1]), 
          .D0(pwm_pulse_level_flag), .A1(n52392), .B1(state_2__N_199_c_1), 
          .C1(time_high_count[2]), .D1(pwm_pulse_level_flag), .CIN(n43926), 
          .COUT(n43927), .S0(time_high_count_15__N_224[1]), .S1(time_high_count_15__N_224[2]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3751_3.INIT0 = 16'hf070;
    defparam add_3751_3.INIT1 = 16'hf070;
    defparam add_3751_3.INJECT1_0 = "NO";
    defparam add_3751_3.INJECT1_1 = "NO";
    CCU2D add_3751_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(time_high_count[0]), .B1(n47131), .C1(state_2__N_199_c_1), 
          .D1(pwm_pulse_level_flag), .COUT(n43926), .S1(time_high_count_15__N_224[0]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3751_1.INIT0 = 16'hF000;
    defparam add_3751_1.INIT1 = 16'hd222;
    defparam add_3751_1.INJECT1_0 = "NO";
    defparam add_3751_1.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut (.A(state[2]), .B(state[1]), .C(state[0]), .D(time_high_count_15__N_224[15]), 
         .Z(time_high_count_15__N_183[15])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_435 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[14]), .Z(time_high_count_15__N_183[14])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_435.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_436 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[13]), .Z(time_high_count_15__N_183[13])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_436.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_437 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[12]), .Z(time_high_count_15__N_183[12])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_437.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_438 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[11]), .Z(time_high_count_15__N_183[11])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_438.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_439 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[10]), .Z(time_high_count_15__N_183[10])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_439.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_440 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[9]), .Z(time_high_count_15__N_183[9])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_440.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_441 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[8]), .Z(time_high_count_15__N_183[8])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_441.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_442 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[7]), .Z(time_high_count_15__N_183[7])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_442.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_443 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[6]), .Z(time_high_count_15__N_183[6])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_443.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_444 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[5]), .Z(time_high_count_15__N_183[5])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_444.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_445 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[4]), .Z(time_high_count_15__N_183[4])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_445.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_446 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[3]), .Z(time_high_count_15__N_183[3])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_446.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_447 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[2]), .Z(time_high_count_15__N_183[2])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_447.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_448 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[1]), .Z(time_high_count_15__N_183[1])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_448.init = 16'h0400;
    PFUMX i40938 (.BLUT(n52516), .ALUT(n52517), .C0(time_high_count[4]), 
          .Z(n52518));
    FD1P3JX time_high_us_i2 (.D(n51098), .SP(us_clk_enable_134), .PD(n30680), 
            .CK(us_clk), .Q(\roll_pwm_pulse_length_us[2] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=52, LSE_RCOL=25, LSE_LLINE=92, LSE_RLINE=98 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i2.GSR = "ENABLED";
    FD1P3JX time_high_us_i3 (.D(n48998), .SP(us_clk_enable_134), .PD(n30680), 
            .CK(us_clk), .Q(\roll_pwm_pulse_length_us[3] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=52, LSE_RCOL=25, LSE_LLINE=92, LSE_RLINE=98 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i3.GSR = "ENABLED";
    FD1P3JX time_high_us_i4 (.D(n52518), .SP(us_clk_enable_134), .PD(n30680), 
            .CK(us_clk), .Q(\roll_pwm_pulse_length_us[4] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=52, LSE_RCOL=25, LSE_LLINE=92, LSE_RLINE=98 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i4.GSR = "ENABLED";
    FD1P3IX time_high_us_i5 (.D(pwm_pulse_length_us_15__N_208[5]), .SP(us_clk_enable_134), 
            .CD(n30680), .CK(us_clk), .Q(\roll_pwm_pulse_length_us[5] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=52, LSE_RCOL=25, LSE_LLINE=92, LSE_RLINE=98 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i5.GSR = "ENABLED";
    FD1P3JX time_high_us_i6 (.D(n3), .SP(us_clk_enable_134), .PD(n30680), 
            .CK(us_clk), .Q(\roll_pwm_pulse_length_us[6] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=52, LSE_RCOL=25, LSE_LLINE=92, LSE_RLINE=98 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i6.GSR = "ENABLED";
    FD1P3JX time_high_us_i7 (.D(n3_adj_5346), .SP(us_clk_enable_134), .PD(n30680), 
            .CK(us_clk), .Q(\roll_pwm_pulse_length_us[7] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=52, LSE_RCOL=25, LSE_LLINE=92, LSE_RLINE=98 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i7.GSR = "ENABLED";
    FD1P3JX time_high_us_i8 (.D(n3_adj_5347), .SP(us_clk_enable_134), .PD(n30680), 
            .CK(us_clk), .Q(\roll_pwm_pulse_length_us[8] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=52, LSE_RCOL=25, LSE_LLINE=92, LSE_RLINE=98 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i8.GSR = "ENABLED";
    FD1P3IX time_high_us_i9 (.D(pwm_pulse_length_us_15__N_208[9]), .SP(us_clk_enable_134), 
            .CD(n30680), .CK(us_clk), .Q(\roll_pwm_pulse_length_us[9] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=52, LSE_RCOL=25, LSE_LLINE=92, LSE_RLINE=98 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i9.GSR = "ENABLED";
    FD1P3IX pwm_pulse_level_flag_46 (.D(n46549), .SP(us_clk_enable_146), 
            .CD(n36401), .CK(us_clk), .Q(pwm_pulse_level_flag)) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=52, LSE_RCOL=25, LSE_LLINE=92, LSE_RLINE=98 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam pwm_pulse_level_flag_46.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module pwm_to_value_U4
//

module pwm_to_value_U4 (latched_roll, us_clk, \roll_pwm_pulse_length_us[2] , 
            \roll_pwm_pulse_length_us[5] , \roll_pwm_pulse_length_us[7] , 
            \roll_pwm_pulse_length_us[6] , \roll_pwm_pulse_length_us[4] , 
            \roll_pwm_pulse_length_us[3] , \roll_pwm_pulse_length_us[8] , 
            n48820, \roll_pwm_pulse_length_us[9] ) /* synthesis syn_module_defined=1 */ ;
    output [7:0]latched_roll;
    input us_clk;
    input \roll_pwm_pulse_length_us[2] ;
    input \roll_pwm_pulse_length_us[5] ;
    input \roll_pwm_pulse_length_us[7] ;
    input \roll_pwm_pulse_length_us[6] ;
    input \roll_pwm_pulse_length_us[4] ;
    input \roll_pwm_pulse_length_us[3] ;
    input \roll_pwm_pulse_length_us[8] ;
    output n48820;
    input \roll_pwm_pulse_length_us[9] ;
    
    wire us_clk /* synthesis SET_AS_NETWORK=us_clk, is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(221[10:16])
    
    wire n52385;
    wire [15:0]value_out_7__N_154;
    
    wire n52266, n52226;
    
    FD1S3AX adjusted_value_i0 (.D(\roll_pwm_pulse_length_us[2] ), .CK(us_clk), 
            .Q(latched_roll[0])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=100, LSE_RLINE=105 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i0.GSR = "DISABLED";
    LUT4 i7404_2_lut_3_lut_4_lut (.A(\roll_pwm_pulse_length_us[5] ), .B(n52385), 
         .C(\roll_pwm_pulse_length_us[7] ), .D(\roll_pwm_pulse_length_us[6] ), 
         .Z(value_out_7__N_154[7])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;
    defparam i7404_2_lut_3_lut_4_lut.init = 16'h78f0;
    FD1S3AX adjusted_value_i7 (.D(value_out_7__N_154[9]), .CK(us_clk), .Q(latched_roll[7])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=100, LSE_RLINE=105 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i7.GSR = "DISABLED";
    FD1S3AX adjusted_value_i6 (.D(value_out_7__N_154[8]), .CK(us_clk), .Q(latched_roll[6])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=100, LSE_RLINE=105 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i6.GSR = "DISABLED";
    FD1S3AX adjusted_value_i5 (.D(value_out_7__N_154[7]), .CK(us_clk), .Q(latched_roll[5])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=100, LSE_RLINE=105 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i5.GSR = "DISABLED";
    FD1S3AX adjusted_value_i4 (.D(value_out_7__N_154[6]), .CK(us_clk), .Q(latched_roll[4])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=100, LSE_RLINE=105 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i4.GSR = "DISABLED";
    FD1S3AX adjusted_value_i3 (.D(value_out_7__N_154[5]), .CK(us_clk), .Q(latched_roll[3])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=100, LSE_RLINE=105 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i3.GSR = "DISABLED";
    FD1S3AX adjusted_value_i2 (.D(value_out_7__N_154[4]), .CK(us_clk), .Q(latched_roll[2])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=100, LSE_RLINE=105 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i2.GSR = "DISABLED";
    FD1S3AX adjusted_value_i1 (.D(value_out_7__N_154[3]), .CK(us_clk), .Q(latched_roll[1])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=100, LSE_RLINE=105 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i1.GSR = "DISABLED";
    LUT4 i7387_2_lut_rep_449 (.A(\roll_pwm_pulse_length_us[4] ), .B(\roll_pwm_pulse_length_us[3] ), 
         .Z(n52385)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i7387_2_lut_rep_449.init = 16'heeee;
    LUT4 i7392_2_lut_rep_330_3_lut (.A(\roll_pwm_pulse_length_us[4] ), .B(\roll_pwm_pulse_length_us[3] ), 
         .C(\roll_pwm_pulse_length_us[5] ), .Z(n52266)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i7392_2_lut_rep_330_3_lut.init = 16'he0e0;
    LUT4 i7390_2_lut_3_lut (.A(\roll_pwm_pulse_length_us[4] ), .B(\roll_pwm_pulse_length_us[3] ), 
         .C(\roll_pwm_pulse_length_us[5] ), .Z(value_out_7__N_154[5])) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B !(C)))) */ ;
    defparam i7390_2_lut_3_lut.init = 16'h1e1e;
    LUT4 i7399_2_lut_rep_290_3_lut_4_lut (.A(\roll_pwm_pulse_length_us[4] ), 
         .B(\roll_pwm_pulse_length_us[3] ), .C(\roll_pwm_pulse_length_us[6] ), 
         .D(\roll_pwm_pulse_length_us[5] ), .Z(n52226)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;
    defparam i7399_2_lut_rep_290_3_lut_4_lut.init = 16'he000;
    LUT4 i7397_2_lut_3_lut_4_lut (.A(\roll_pwm_pulse_length_us[4] ), .B(\roll_pwm_pulse_length_us[3] ), 
         .C(\roll_pwm_pulse_length_us[6] ), .D(\roll_pwm_pulse_length_us[5] ), 
         .Z(value_out_7__N_154[6])) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B !(C)))) */ ;
    defparam i7397_2_lut_3_lut_4_lut.init = 16'h1ef0;
    LUT4 i1_2_lut (.A(\roll_pwm_pulse_length_us[4] ), .B(\roll_pwm_pulse_length_us[3] ), 
         .Z(value_out_7__N_154[4])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i1_2_lut.init = 16'h9999;
    LUT4 i7380_1_lut (.A(\roll_pwm_pulse_length_us[3] ), .Z(value_out_7__N_154[3])) /* synthesis lut_function=(!(A)) */ ;
    defparam i7380_1_lut.init = 16'h5555;
    LUT4 i7411_2_lut_3_lut_4_lut (.A(\roll_pwm_pulse_length_us[6] ), .B(n52266), 
         .C(\roll_pwm_pulse_length_us[8] ), .D(\roll_pwm_pulse_length_us[7] ), 
         .Z(value_out_7__N_154[8])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;
    defparam i7411_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i2_3_lut (.A(latched_roll[2]), .B(latched_roll[1]), .C(latched_roll[3]), 
         .Z(n48820)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i2_3_lut.init = 16'h1010;
    LUT4 i7418_3_lut_4_lut (.A(\roll_pwm_pulse_length_us[7] ), .B(n52226), 
         .C(\roll_pwm_pulse_length_us[8] ), .D(\roll_pwm_pulse_length_us[9] ), 
         .Z(value_out_7__N_154[9])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;
    defparam i7418_3_lut_4_lut.init = 16'h7f80;
    
endmodule
//
// Verilog Description of module pwm_reader_U5
//

module pwm_reader_U5 (state_2__N_199_c_1, us_clk, GND_net, \pitch_pwm_pulse_length_us[2] , 
            \pitch_pwm_pulse_length_us[3] , \pitch_pwm_pulse_length_us[4] , 
            \pitch_pwm_pulse_length_us[5] , \pitch_pwm_pulse_length_us[6] , 
            \pitch_pwm_pulse_length_us[7] , \pitch_pwm_pulse_length_us[8] , 
            \pitch_pwm_pulse_length_us[9] ) /* synthesis syn_module_defined=1 */ ;
    input state_2__N_199_c_1;
    input us_clk;
    input GND_net;
    output \pitch_pwm_pulse_length_us[2] ;
    output \pitch_pwm_pulse_length_us[3] ;
    output \pitch_pwm_pulse_length_us[4] ;
    output \pitch_pwm_pulse_length_us[5] ;
    output \pitch_pwm_pulse_length_us[6] ;
    output \pitch_pwm_pulse_length_us[7] ;
    output \pitch_pwm_pulse_length_us[8] ;
    output \pitch_pwm_pulse_length_us[9] ;
    
    wire us_clk /* synthesis SET_AS_NETWORK=us_clk, is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(221[10:16])
    wire [2:0]state;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(54[15:20])
    
    wire us_clk_enable_145;
    wire [15:0]time_high_count;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(57[16:31])
    
    wire us_clk_enable_18;
    wire [15:0]time_high_count_15__N_183;
    wire [2:0]state_2__N_180;
    
    wire n46783, us_clk_enable_20, n4, pwm_pulse_level_flag, n48982, 
        n18, n16, n16_adj_5343, n16_adj_5344, n47338, n52220, n51056, 
        n51057, n106;
    wire [15:0]pwm_pulse_length_us_15__N_208;
    
    wire n52382, n47133;
    wire [15:0]time_high_count_15__N_224;
    
    wire n48070, n30659, us_clk_enable_143, n49066, n47785, n12, 
        n5, n6, n6_adj_5345, n37360, n3, n48817, n36407, n46515, 
        n43909, n43908, n43907, n43906, n43905, n43904, n43903, 
        n43902;
    
    LUT4 i20_4_lut_3_lut_4_lut (.A(state[1]), .B(state_2__N_199_c_1), .C(state[0]), 
         .D(state[2]), .Z(us_clk_enable_145)) /* synthesis lut_function=(A (B ((D)+!C)+!B (D))+!A !(D)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(74[13] 161[20])
    defparam i20_4_lut_3_lut_4_lut.init = 16'haa5d;
    FD1P3AX time_high_count_i0 (.D(time_high_count_15__N_183[0]), .SP(us_clk_enable_18), 
            .CK(us_clk), .Q(time_high_count[0])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=53, LSE_RCOL=25, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i0.GSR = "ENABLED";
    FD1S3AX state_i0 (.D(state_2__N_180[0]), .CK(us_clk), .Q(state[0])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=14, LSE_LCOL=53, LSE_RCOL=25, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam state_i0.GSR = "ENABLED";
    FD1S3IX state_i2 (.D(n46783), .CK(us_clk), .CD(state[2]), .Q(state[2])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=14, LSE_LCOL=53, LSE_RCOL=25, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam state_i2.GSR = "ENABLED";
    FD1S3AX state_i1 (.D(state_2__N_180[1]), .CK(us_clk), .Q(state[1])) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=14, LSE_LCOL=53, LSE_RCOL=25, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam state_i1.GSR = "ENABLED";
    FD1P3AX time_high_count_i15 (.D(time_high_count_15__N_183[15]), .SP(us_clk_enable_18), 
            .CK(us_clk), .Q(time_high_count[15])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=53, LSE_RCOL=25, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i15.GSR = "ENABLED";
    FD1P3AX time_high_count_i14 (.D(time_high_count_15__N_183[14]), .SP(us_clk_enable_18), 
            .CK(us_clk), .Q(time_high_count[14])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=53, LSE_RCOL=25, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i14.GSR = "ENABLED";
    FD1P3AX time_high_count_i13 (.D(time_high_count_15__N_183[13]), .SP(us_clk_enable_18), 
            .CK(us_clk), .Q(time_high_count[13])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=53, LSE_RCOL=25, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i13.GSR = "ENABLED";
    FD1P3AX time_high_count_i12 (.D(time_high_count_15__N_183[12]), .SP(us_clk_enable_18), 
            .CK(us_clk), .Q(time_high_count[12])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=53, LSE_RCOL=25, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i12.GSR = "ENABLED";
    FD1P3AX time_high_count_i11 (.D(time_high_count_15__N_183[11]), .SP(us_clk_enable_18), 
            .CK(us_clk), .Q(time_high_count[11])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=53, LSE_RCOL=25, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i11.GSR = "ENABLED";
    FD1P3AX time_high_count_i10 (.D(time_high_count_15__N_183[10]), .SP(us_clk_enable_18), 
            .CK(us_clk), .Q(time_high_count[10])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=53, LSE_RCOL=25, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i10.GSR = "ENABLED";
    FD1P3AX time_high_count_i9 (.D(time_high_count_15__N_183[9]), .SP(us_clk_enable_18), 
            .CK(us_clk), .Q(time_high_count[9])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=53, LSE_RCOL=25, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i9.GSR = "ENABLED";
    FD1P3AX time_high_count_i8 (.D(time_high_count_15__N_183[8]), .SP(us_clk_enable_18), 
            .CK(us_clk), .Q(time_high_count[8])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=53, LSE_RCOL=25, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i8.GSR = "ENABLED";
    FD1P3AX time_high_count_i7 (.D(time_high_count_15__N_183[7]), .SP(us_clk_enable_18), 
            .CK(us_clk), .Q(time_high_count[7])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=53, LSE_RCOL=25, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i7.GSR = "ENABLED";
    FD1P3AX time_high_count_i6 (.D(time_high_count_15__N_183[6]), .SP(us_clk_enable_18), 
            .CK(us_clk), .Q(time_high_count[6])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=53, LSE_RCOL=25, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i6.GSR = "ENABLED";
    FD1P3AX time_high_count_i5 (.D(time_high_count_15__N_183[5]), .SP(us_clk_enable_18), 
            .CK(us_clk), .Q(time_high_count[5])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=53, LSE_RCOL=25, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i5.GSR = "ENABLED";
    FD1P3AX time_high_count_i4 (.D(time_high_count_15__N_183[4]), .SP(us_clk_enable_18), 
            .CK(us_clk), .Q(time_high_count[4])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=53, LSE_RCOL=25, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i4.GSR = "ENABLED";
    FD1P3AX time_high_count_i3 (.D(time_high_count_15__N_183[3]), .SP(us_clk_enable_18), 
            .CK(us_clk), .Q(time_high_count[3])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=53, LSE_RCOL=25, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i3.GSR = "ENABLED";
    FD1P3AX time_high_count_i2 (.D(time_high_count_15__N_183[2]), .SP(us_clk_enable_20), 
            .CK(us_clk), .Q(time_high_count[2])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=53, LSE_RCOL=25, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i2.GSR = "ENABLED";
    FD1P3AX time_high_count_i1 (.D(time_high_count_15__N_183[1]), .SP(us_clk_enable_20), 
            .CK(us_clk), .Q(time_high_count[1])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=53, LSE_RCOL=25, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_count_i1.GSR = "ENABLED";
    LUT4 i2_4_lut (.A(state[0]), .B(state_2__N_199_c_1), .C(state[1]), 
         .D(n4), .Z(us_clk_enable_18)) /* synthesis lut_function=((B (C)+!B (C+!(D)))+!A) */ ;
    defparam i2_4_lut.init = 16'hf5f7;
    LUT4 i1_2_lut (.A(state[2]), .B(pwm_pulse_level_flag), .Z(n4)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i39604_3_lut_4_lut (.A(n48982), .B(n18), .C(time_high_count[6]), 
         .D(state[1]), .Z(n16)) /* synthesis lut_function=(A (D)+!A (B (C (D))+!B (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(74[13] 161[20])
    defparam i39604_3_lut_4_lut.init = 16'hfb00;
    LUT4 i39614_3_lut_4_lut (.A(n48982), .B(n18), .C(time_high_count[7]), 
         .D(state[1]), .Z(n16_adj_5343)) /* synthesis lut_function=(A (D)+!A (B (C (D))+!B (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(74[13] 161[20])
    defparam i39614_3_lut_4_lut.init = 16'hfb00;
    LUT4 i39619_3_lut_4_lut (.A(n48982), .B(n18), .C(time_high_count[8]), 
         .D(state[1]), .Z(n16_adj_5344)) /* synthesis lut_function=(A (D)+!A (B (C (D))+!B (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(74[13] 161[20])
    defparam i39619_3_lut_4_lut.init = 16'hfb00;
    LUT4 i1_2_lut_rep_284 (.A(n47338), .B(n18), .Z(n52220)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_284.init = 16'heeee;
    LUT4 state_1__bdd_3_lut (.A(state[1]), .B(state[0]), .C(state_2__N_199_c_1), 
         .Z(n51056)) /* synthesis lut_function=(!(A+!((C)+!B))) */ ;
    defparam state_1__bdd_3_lut.init = 16'h5151;
    LUT4 state_1__bdd_4_lut (.A(state[1]), .B(pwm_pulse_level_flag), .C(state[0]), 
         .D(state_2__N_199_c_1), .Z(n51057)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A (((D)+!C)+!B))) */ ;
    defparam state_1__bdd_4_lut.init = 16'h0840;
    LUT4 i25871_3_lut_4_lut (.A(n47338), .B(n18), .C(n106), .D(time_high_count[5]), 
         .Z(pwm_pulse_length_us_15__N_208[5])) /* synthesis lut_function=(!(A (C+!(D))+!A (B (C+!(D))))) */ ;
    defparam i25871_3_lut_4_lut.init = 16'h1f11;
    LUT4 state_0__bdd_4_lut (.A(state[0]), .B(state[2]), .C(state[1]), 
         .D(state_2__N_199_c_1), .Z(state_2__N_180[0])) /* synthesis lut_function=(!(A (B (C+(D)))+!A (B+(C (D))))) */ ;
    defparam state_0__bdd_4_lut.init = 16'h233b;
    LUT4 pwm_pulse_level_flag_I_0_55_1_lut_rep_446 (.A(pwm_pulse_level_flag), 
         .Z(n52382)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[46:74])
    defparam pwm_pulse_level_flag_I_0_55_1_lut_rep_446.init = 16'h5555;
    LUT4 i1_2_lut_2_lut (.A(pwm_pulse_level_flag), .B(state_2__N_199_c_1), 
         .Z(n47133)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[46:74])
    defparam i1_2_lut_2_lut.init = 16'h4444;
    LUT4 i21_4_lut (.A(state_2__N_199_c_1), .B(pwm_pulse_level_flag), .C(state[1]), 
         .D(state[0]), .Z(n46783)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A ((D)+!C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(74[13] 161[20])
    defparam i21_4_lut.init = 16'h0a70;
    LUT4 i1_2_lut_4_lut (.A(state[2]), .B(state[1]), .C(state[0]), .D(time_high_count_15__N_224[15]), 
         .Z(time_high_count_15__N_183[15])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_406 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[14]), .Z(time_high_count_15__N_183[14])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_406.init = 16'h0400;
    LUT4 i39954_4_lut (.A(pwm_pulse_level_flag), .B(n48070), .C(state_2__N_199_c_1), 
         .D(state[2]), .Z(us_clk_enable_20)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))))) */ ;
    defparam i39954_4_lut.init = 16'h3337;
    LUT4 i1_2_lut_4_lut_adj_407 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[13]), .Z(time_high_count_15__N_183[13])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_407.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_408 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[12]), .Z(time_high_count_15__N_183[12])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_408.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_409 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[11]), .Z(time_high_count_15__N_183[11])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_409.init = 16'h0400;
    LUT4 i1_2_lut_adj_410 (.A(state[1]), .B(state[0]), .Z(n48070)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_adj_410.init = 16'h4444;
    LUT4 i1_2_lut_4_lut_adj_411 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[10]), .Z(time_high_count_15__N_183[10])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_411.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_412 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[9]), .Z(time_high_count_15__N_183[9])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_412.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_413 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[8]), .Z(time_high_count_15__N_183[8])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_413.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_414 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[7]), .Z(time_high_count_15__N_183[7])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_414.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_415 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[6]), .Z(time_high_count_15__N_183[6])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_415.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_416 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[5]), .Z(time_high_count_15__N_183[5])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_416.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_417 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[4]), .Z(time_high_count_15__N_183[4])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_417.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_418 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[3]), .Z(time_high_count_15__N_183[3])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_418.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_419 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[2]), .Z(time_high_count_15__N_183[2])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_419.init = 16'h0400;
    LUT4 i1_2_lut_4_lut_adj_420 (.A(state[2]), .B(state[1]), .C(state[0]), 
         .D(time_high_count_15__N_224[1]), .Z(time_high_count_15__N_183[1])) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i1_2_lut_4_lut_adj_420.init = 16'h0400;
    LUT4 i2_3_lut_4_lut (.A(state[1]), .B(state[2]), .C(time_high_count_15__N_224[0]), 
         .D(state[0]), .Z(time_high_count_15__N_183[0])) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i2_3_lut_4_lut.init = 16'h0020;
    LUT4 i19995_2_lut_4_lut_3_lut (.A(state[1]), .B(state[2]), .C(state[0]), 
         .Z(n30659)) /* synthesis lut_function=(A (B)+!A !(B+(C))) */ ;
    defparam i19995_2_lut_4_lut_3_lut.init = 16'h8989;
    LUT4 i39410_3_lut_rep_413 (.A(state[0]), .B(state[1]), .C(state[2]), 
         .Z(us_clk_enable_143)) /* synthesis lut_function=(A (B)+!A (B (C)+!B !(C))) */ ;
    defparam i39410_3_lut_rep_413.init = 16'hc9c9;
    PFUMX i40209 (.BLUT(n51057), .ALUT(n51056), .C0(state[2]), .Z(state_2__N_180[1]));
    LUT4 i3_4_lut (.A(state[1]), .B(n106), .C(time_high_count[2]), .D(n52220), 
         .Z(n49066)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i3_4_lut.init = 16'h2000;
    LUT4 i1_4_lut (.A(time_high_count[10]), .B(n47338), .C(n47785), .D(n12), 
         .Z(n106)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;
    defparam i1_4_lut.init = 16'heccc;
    LUT4 i7211_4_lut (.A(n5), .B(time_high_count[5]), .C(time_high_count[4]), 
         .D(n6), .Z(n12)) /* synthesis lut_function=(A (B+(C))+!A (B+(C (D)))) */ ;
    defparam i7211_4_lut.init = 16'hfcec;
    LUT4 i1_2_lut_adj_421 (.A(time_high_count[0]), .B(time_high_count[3]), 
         .Z(n5)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_421.init = 16'heeee;
    LUT4 i2_2_lut (.A(time_high_count[1]), .B(time_high_count[2]), .Z(n6)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i4_4_lut (.A(time_high_count[13]), .B(time_high_count[11]), .C(time_high_count[15]), 
         .D(n6_adj_5345), .Z(n47338)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i4_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_422 (.A(time_high_count[10]), .B(time_high_count[5]), 
         .C(n47785), .D(n37360), .Z(n18)) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(74[13] 161[20])
    defparam i1_4_lut_adj_422.init = 16'heaaa;
    LUT4 i26711_2_lut (.A(time_high_count[3]), .B(time_high_count[4]), .Z(n37360)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i26711_2_lut.init = 16'heeee;
    LUT4 i3_4_lut_adj_423 (.A(time_high_count[9]), .B(time_high_count[6]), 
         .C(time_high_count[8]), .D(time_high_count[7]), .Z(n47785)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i3_4_lut_adj_423.init = 16'h8000;
    LUT4 i1_2_lut_adj_424 (.A(time_high_count[12]), .B(time_high_count[14]), 
         .Z(n6_adj_5345)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_424.init = 16'heeee;
    LUT4 i26911_4_lut (.A(time_high_count[3]), .B(state[1]), .C(n52220), 
         .D(n106), .Z(n3)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A ((C)+!B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(74[13] 161[20])
    defparam i26911_4_lut.init = 16'h0c8c;
    LUT4 i2_4_lut_adj_425 (.A(n52220), .B(state[1]), .C(time_high_count[4]), 
         .D(n106), .Z(n48817)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(74[13] 161[20])
    defparam i2_4_lut_adj_425.init = 16'h8880;
    LUT4 i4_4_lut_adj_426 (.A(time_high_count[13]), .B(time_high_count[15]), 
         .C(time_high_count[11]), .D(n6_adj_5345), .Z(n48982)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i4_4_lut_adj_426.init = 16'hfffe;
    LUT4 i39901_3_lut (.A(time_high_count[9]), .B(n48982), .C(time_high_count[10]), 
         .Z(pwm_pulse_length_us_15__N_208[9])) /* synthesis lut_function=(A+(B+!(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(135[30] 138[65])
    defparam i39901_3_lut.init = 16'hefef;
    LUT4 i25786_2_lut (.A(state[2]), .B(state[1]), .Z(n36407)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam i25786_2_lut.init = 16'h8888;
    LUT4 i1_4_lut_adj_427 (.A(pwm_pulse_level_flag), .B(state[1]), .C(state_2__N_199_c_1), 
         .D(state[0]), .Z(n46515)) /* synthesis lut_function=(A (B+(C (D)))+!A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(74[13] 161[20])
    defparam i1_4_lut_adj_427.init = 16'heccc;
    CCU2D add_3755_17 (.A0(n52382), .B0(state_2__N_199_c_1), .C0(time_high_count[15]), 
          .D0(pwm_pulse_level_flag), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43909), .S0(time_high_count_15__N_224[15]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3755_17.INIT0 = 16'hf070;
    defparam add_3755_17.INIT1 = 16'h0000;
    defparam add_3755_17.INJECT1_0 = "NO";
    defparam add_3755_17.INJECT1_1 = "NO";
    CCU2D add_3755_15 (.A0(n52382), .B0(state_2__N_199_c_1), .C0(time_high_count[13]), 
          .D0(pwm_pulse_level_flag), .A1(n52382), .B1(state_2__N_199_c_1), 
          .C1(time_high_count[14]), .D1(pwm_pulse_level_flag), .CIN(n43908), 
          .COUT(n43909), .S0(time_high_count_15__N_224[13]), .S1(time_high_count_15__N_224[14]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3755_15.INIT0 = 16'hf070;
    defparam add_3755_15.INIT1 = 16'hf070;
    defparam add_3755_15.INJECT1_0 = "NO";
    defparam add_3755_15.INJECT1_1 = "NO";
    CCU2D add_3755_13 (.A0(n52382), .B0(state_2__N_199_c_1), .C0(time_high_count[11]), 
          .D0(pwm_pulse_level_flag), .A1(n52382), .B1(state_2__N_199_c_1), 
          .C1(time_high_count[12]), .D1(pwm_pulse_level_flag), .CIN(n43907), 
          .COUT(n43908), .S0(time_high_count_15__N_224[11]), .S1(time_high_count_15__N_224[12]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3755_13.INIT0 = 16'hf070;
    defparam add_3755_13.INIT1 = 16'hf070;
    defparam add_3755_13.INJECT1_0 = "NO";
    defparam add_3755_13.INJECT1_1 = "NO";
    CCU2D add_3755_11 (.A0(n52382), .B0(state_2__N_199_c_1), .C0(time_high_count[9]), 
          .D0(pwm_pulse_level_flag), .A1(n52382), .B1(state_2__N_199_c_1), 
          .C1(time_high_count[10]), .D1(pwm_pulse_level_flag), .CIN(n43906), 
          .COUT(n43907), .S0(time_high_count_15__N_224[9]), .S1(time_high_count_15__N_224[10]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3755_11.INIT0 = 16'hf070;
    defparam add_3755_11.INIT1 = 16'hf070;
    defparam add_3755_11.INJECT1_0 = "NO";
    defparam add_3755_11.INJECT1_1 = "NO";
    CCU2D add_3755_9 (.A0(n52382), .B0(state_2__N_199_c_1), .C0(time_high_count[7]), 
          .D0(pwm_pulse_level_flag), .A1(n52382), .B1(state_2__N_199_c_1), 
          .C1(time_high_count[8]), .D1(pwm_pulse_level_flag), .CIN(n43905), 
          .COUT(n43906), .S0(time_high_count_15__N_224[7]), .S1(time_high_count_15__N_224[8]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3755_9.INIT0 = 16'hf070;
    defparam add_3755_9.INIT1 = 16'hf070;
    defparam add_3755_9.INJECT1_0 = "NO";
    defparam add_3755_9.INJECT1_1 = "NO";
    CCU2D add_3755_7 (.A0(n52382), .B0(state_2__N_199_c_1), .C0(time_high_count[5]), 
          .D0(pwm_pulse_level_flag), .A1(n52382), .B1(state_2__N_199_c_1), 
          .C1(time_high_count[6]), .D1(pwm_pulse_level_flag), .CIN(n43904), 
          .COUT(n43905), .S0(time_high_count_15__N_224[5]), .S1(time_high_count_15__N_224[6]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3755_7.INIT0 = 16'hf070;
    defparam add_3755_7.INIT1 = 16'hf070;
    defparam add_3755_7.INJECT1_0 = "NO";
    defparam add_3755_7.INJECT1_1 = "NO";
    CCU2D add_3755_5 (.A0(n52382), .B0(state_2__N_199_c_1), .C0(time_high_count[3]), 
          .D0(pwm_pulse_level_flag), .A1(n52382), .B1(state_2__N_199_c_1), 
          .C1(time_high_count[4]), .D1(pwm_pulse_level_flag), .CIN(n43903), 
          .COUT(n43904), .S0(time_high_count_15__N_224[3]), .S1(time_high_count_15__N_224[4]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3755_5.INIT0 = 16'hf070;
    defparam add_3755_5.INIT1 = 16'hf070;
    defparam add_3755_5.INJECT1_0 = "NO";
    defparam add_3755_5.INJECT1_1 = "NO";
    CCU2D add_3755_3 (.A0(n52382), .B0(state_2__N_199_c_1), .C0(time_high_count[1]), 
          .D0(pwm_pulse_level_flag), .A1(n52382), .B1(state_2__N_199_c_1), 
          .C1(time_high_count[2]), .D1(pwm_pulse_level_flag), .CIN(n43902), 
          .COUT(n43903), .S0(time_high_count_15__N_224[1]), .S1(time_high_count_15__N_224[2]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3755_3.INIT0 = 16'hf070;
    defparam add_3755_3.INIT1 = 16'hf070;
    defparam add_3755_3.INJECT1_0 = "NO";
    defparam add_3755_3.INJECT1_1 = "NO";
    CCU2D add_3755_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(time_high_count[0]), .B1(n47133), .C1(state_2__N_199_c_1), 
          .D1(pwm_pulse_level_flag), .COUT(n43902), .S1(time_high_count_15__N_224[0]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(115[26] 125[24])
    defparam add_3755_1.INIT0 = 16'hF000;
    defparam add_3755_1.INIT1 = 16'hd222;
    defparam add_3755_1.INJECT1_0 = "NO";
    defparam add_3755_1.INJECT1_1 = "NO";
    FD1P3JX time_high_us_i2 (.D(n49066), .SP(us_clk_enable_143), .PD(n30659), 
            .CK(us_clk), .Q(\pitch_pwm_pulse_length_us[2] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=53, LSE_RCOL=25, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i2.GSR = "ENABLED";
    FD1P3JX time_high_us_i3 (.D(n3), .SP(us_clk_enable_143), .PD(n30659), 
            .CK(us_clk), .Q(\pitch_pwm_pulse_length_us[3] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=53, LSE_RCOL=25, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i3.GSR = "ENABLED";
    FD1P3JX time_high_us_i4 (.D(n48817), .SP(us_clk_enable_143), .PD(n30659), 
            .CK(us_clk), .Q(\pitch_pwm_pulse_length_us[4] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=53, LSE_RCOL=25, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i4.GSR = "ENABLED";
    FD1P3IX time_high_us_i5 (.D(pwm_pulse_length_us_15__N_208[5]), .SP(us_clk_enable_143), 
            .CD(n30659), .CK(us_clk), .Q(\pitch_pwm_pulse_length_us[5] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=53, LSE_RCOL=25, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i5.GSR = "ENABLED";
    FD1P3JX time_high_us_i6 (.D(n16), .SP(us_clk_enable_143), .PD(n30659), 
            .CK(us_clk), .Q(\pitch_pwm_pulse_length_us[6] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=53, LSE_RCOL=25, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i6.GSR = "ENABLED";
    FD1P3JX time_high_us_i7 (.D(n16_adj_5343), .SP(us_clk_enable_143), .PD(n30659), 
            .CK(us_clk), .Q(\pitch_pwm_pulse_length_us[7] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=53, LSE_RCOL=25, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i7.GSR = "ENABLED";
    FD1P3JX time_high_us_i8 (.D(n16_adj_5344), .SP(us_clk_enable_143), .PD(n30659), 
            .CK(us_clk), .Q(\pitch_pwm_pulse_length_us[8] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=53, LSE_RCOL=25, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i8.GSR = "ENABLED";
    FD1P3IX time_high_us_i9 (.D(pwm_pulse_length_us_15__N_208[9]), .SP(us_clk_enable_143), 
            .CD(n30659), .CK(us_clk), .Q(\pitch_pwm_pulse_length_us[9] )) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=53, LSE_RCOL=25, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam time_high_us_i9.GSR = "ENABLED";
    FD1P3IX pwm_pulse_level_flag_46 (.D(n46515), .SP(us_clk_enable_145), 
            .CD(n36407), .CK(us_clk), .Q(pwm_pulse_level_flag)) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=53, LSE_RCOL=25, LSE_LLINE=108, LSE_RLINE=114 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_reader.v(73[14] 162[12])
    defparam pwm_pulse_level_flag_46.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module pwm_to_value_U6
//

module pwm_to_value_U6 (\latched_roll[2] , \latched_roll[3] , \latched_roll[1] , 
            n1406, latched_pitch, us_clk, \pitch_pwm_pulse_length_us[2] , 
            n52328, \tx_byte_index[0] , n52095, n27, \tx_byte_index[1] , 
            \tx_word_index[1] , n36649, n34665, \pitch_pwm_pulse_length_us[5] , 
            \pitch_pwm_pulse_length_us[7] , \pitch_pwm_pulse_length_us[6] , 
            \pitch_pwm_pulse_length_us[4] , \pitch_pwm_pulse_length_us[3] , 
            n51272, n51271, n51273, \latched_roll[0] , n51202, n51159, 
            \swa_swb_val[0] , \swa_swb_val[1] , \swa_swb_val[2] , \swa_swb_val[3] , 
            n51201, n34692, n36752, \pitch_pwm_pulse_length_us[8] , 
            n34690, \pitch_pwm_pulse_length_us[9] ) /* synthesis syn_module_defined=1 */ ;
    input \latched_roll[2] ;
    input \latched_roll[3] ;
    input \latched_roll[1] ;
    output n1406;
    output [7:0]latched_pitch;
    input us_clk;
    input \pitch_pwm_pulse_length_us[2] ;
    input n52328;
    input \tx_byte_index[0] ;
    output n52095;
    output n27;
    input \tx_byte_index[1] ;
    input \tx_word_index[1] ;
    input n36649;
    output n34665;
    input \pitch_pwm_pulse_length_us[5] ;
    input \pitch_pwm_pulse_length_us[7] ;
    input \pitch_pwm_pulse_length_us[6] ;
    input \pitch_pwm_pulse_length_us[4] ;
    input \pitch_pwm_pulse_length_us[3] ;
    input n51272;
    input n51271;
    output n51273;
    input \latched_roll[0] ;
    output n51202;
    output n51159;
    input \swa_swb_val[0] ;
    input \swa_swb_val[1] ;
    input \swa_swb_val[2] ;
    input \swa_swb_val[3] ;
    output n51201;
    output n34692;
    output n36752;
    input \pitch_pwm_pulse_length_us[8] ;
    output n34690;
    input \pitch_pwm_pulse_length_us[9] ;
    
    wire us_clk /* synthesis SET_AS_NETWORK=us_clk, is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(221[10:16])
    wire [15:0]value_out_7__N_154;
    
    wire n34679, n52427, n13, n52284, n52236;
    
    LUT4 i1_3_lut (.A(\latched_roll[2] ), .B(\latched_roll[3] ), .C(\latched_roll[1] ), 
         .Z(n1406)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/angle_controller.v(84[74:86])
    defparam i1_3_lut.init = 16'hc8c8;
    FD1S3AX adjusted_value_i0 (.D(\pitch_pwm_pulse_length_us[2] ), .CK(us_clk), 
            .Q(latched_pitch[0])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=116, LSE_RLINE=121 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i0.GSR = "DISABLED";
    FD1S3AX adjusted_value_i7 (.D(value_out_7__N_154[9]), .CK(us_clk), .Q(latched_pitch[7])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=116, LSE_RLINE=121 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i7.GSR = "DISABLED";
    FD1S3AX adjusted_value_i6 (.D(value_out_7__N_154[8]), .CK(us_clk), .Q(latched_pitch[6])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=116, LSE_RLINE=121 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i6.GSR = "DISABLED";
    FD1S3AX adjusted_value_i5 (.D(value_out_7__N_154[7]), .CK(us_clk), .Q(latched_pitch[5])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=116, LSE_RLINE=121 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i5.GSR = "DISABLED";
    FD1S3AX adjusted_value_i4 (.D(value_out_7__N_154[6]), .CK(us_clk), .Q(latched_pitch[4])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=116, LSE_RLINE=121 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i4.GSR = "DISABLED";
    FD1S3AX adjusted_value_i3 (.D(value_out_7__N_154[5]), .CK(us_clk), .Q(latched_pitch[3])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=116, LSE_RLINE=121 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i3.GSR = "DISABLED";
    FD1S3AX adjusted_value_i2 (.D(value_out_7__N_154[4]), .CK(us_clk), .Q(latched_pitch[2])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=116, LSE_RLINE=121 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i2.GSR = "DISABLED";
    FD1S3AX adjusted_value_i1 (.D(value_out_7__N_154[3]), .CK(us_clk), .Q(latched_pitch[1])) /* synthesis LSE_LINE_FILE_ID=14, LSE_LCOL=18, LSE_RCOL=25, LSE_LLINE=116, LSE_RLINE=121 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam adjusted_value_i1.GSR = "DISABLED";
    LUT4 n34679_bdd_3_lut_4_lut (.A(n52328), .B(latched_pitch[6]), .C(\tx_byte_index[0] ), 
         .D(n34679), .Z(n52095)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B ((D)+!C))) */ ;
    defparam n34679_bdd_3_lut_4_lut.init = 16'hf101;
    LUT4 i24025_4_lut (.A(n27), .B(\tx_byte_index[1] ), .C(\tx_word_index[1] ), 
         .D(n36649), .Z(n34665)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(97[17:30])
    defparam i24025_4_lut.init = 16'hfaca;
    LUT4 i7455_2_lut_3_lut_4_lut (.A(\pitch_pwm_pulse_length_us[5] ), .B(n52427), 
         .C(\pitch_pwm_pulse_length_us[7] ), .D(\pitch_pwm_pulse_length_us[6] ), 
         .Z(value_out_7__N_154[7])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;
    defparam i7455_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i1_2_lut (.A(\pitch_pwm_pulse_length_us[4] ), .B(\pitch_pwm_pulse_length_us[3] ), 
         .Z(value_out_7__N_154[4])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i1_2_lut.init = 16'h9999;
    LUT4 i7431_1_lut (.A(\pitch_pwm_pulse_length_us[3] ), .Z(value_out_7__N_154[3])) /* synthesis lut_function=(!(A)) */ ;
    defparam i7431_1_lut.init = 16'h5555;
    PFUMX i40332 (.BLUT(n51272), .ALUT(n51271), .C0(\tx_word_index[1] ), 
          .Z(n51273));
    LUT4 swa_swb_val_0__bdd_3_lut_4_lut (.A(\latched_roll[0] ), .B(\latched_roll[3] ), 
         .C(\latched_roll[2] ), .D(\latched_roll[1] ), .Z(n51202)) /* synthesis lut_function=(!(A (C)+!A (B (C (D))+!B (C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/angle_controller.v(84[74:86])
    defparam swa_swb_val_0__bdd_3_lut_4_lut.init = 16'h0f4f;
    LUT4 i8_3_lut_3_lut (.A(latched_pitch[3]), .B(latched_pitch[1]), .C(latched_pitch[2]), 
         .Z(n34679)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam i8_3_lut_3_lut.init = 16'h0202;
    LUT4 i1_4_lut_4_lut (.A(latched_pitch[3]), .B(n13), .C(latched_pitch[2]), 
         .D(\tx_byte_index[1] ), .Z(n27)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (C+(D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_to_value.v(33[20] 36[16])
    defparam i1_4_lut_4_lut.init = 16'hffd0;
    LUT4 i1_2_lut_adj_405 (.A(latched_pitch[1]), .B(latched_pitch[0]), .Z(n13)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_405.init = 16'heeee;
    LUT4 latched_roll_2__bdd_4_lut_41079 (.A(\latched_roll[2] ), .B(\latched_roll[1] ), 
         .C(\latched_roll[3] ), .D(\latched_roll[0] ), .Z(n51159)) /* synthesis lut_function=(A (B ((D)+!C)+!B !((D)+!C))+!A (B ((D)+!C))) */ ;
    defparam latched_roll_2__bdd_4_lut_41079.init = 16'hcc2c;
    LUT4 swa_swb_val_0__bdd_4_lut (.A(\swa_swb_val[0] ), .B(\swa_swb_val[1] ), 
         .C(\swa_swb_val[2] ), .D(\swa_swb_val[3] ), .Z(n51201)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B !((D)+!C)))) */ ;
    defparam swa_swb_val_0__bdd_4_lut.init = 16'h1f0f;
    LUT4 i12_2_lut (.A(\latched_roll[0] ), .B(\latched_roll[3] ), .Z(n34692)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/angle_controller.v(84[74:86])
    defparam i12_2_lut.init = 16'h6666;
    LUT4 i26120_4_lut_3_lut (.A(latched_pitch[1]), .B(latched_pitch[0]), 
         .C(latched_pitch[2]), .Z(n36752)) /* synthesis lut_function=(A (B)+!A !(B+!(C))) */ ;
    defparam i26120_4_lut_3_lut.init = 16'h9898;
    LUT4 i7438_2_lut_rep_491 (.A(\pitch_pwm_pulse_length_us[4] ), .B(\pitch_pwm_pulse_length_us[3] ), 
         .Z(n52427)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i7438_2_lut_rep_491.init = 16'heeee;
    LUT4 i7443_2_lut_rep_348_3_lut (.A(\pitch_pwm_pulse_length_us[4] ), .B(\pitch_pwm_pulse_length_us[3] ), 
         .C(\pitch_pwm_pulse_length_us[5] ), .Z(n52284)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i7443_2_lut_rep_348_3_lut.init = 16'he0e0;
    LUT4 i7441_2_lut_3_lut (.A(\pitch_pwm_pulse_length_us[4] ), .B(\pitch_pwm_pulse_length_us[3] ), 
         .C(\pitch_pwm_pulse_length_us[5] ), .Z(value_out_7__N_154[5])) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B !(C)))) */ ;
    defparam i7441_2_lut_3_lut.init = 16'h1e1e;
    LUT4 i7450_2_lut_rep_300_3_lut_4_lut (.A(\pitch_pwm_pulse_length_us[4] ), 
         .B(\pitch_pwm_pulse_length_us[3] ), .C(\pitch_pwm_pulse_length_us[6] ), 
         .D(\pitch_pwm_pulse_length_us[5] ), .Z(n52236)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;
    defparam i7450_2_lut_rep_300_3_lut_4_lut.init = 16'he000;
    LUT4 i7448_2_lut_3_lut_4_lut (.A(\pitch_pwm_pulse_length_us[4] ), .B(\pitch_pwm_pulse_length_us[3] ), 
         .C(\pitch_pwm_pulse_length_us[6] ), .D(\pitch_pwm_pulse_length_us[5] ), 
         .Z(value_out_7__N_154[6])) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B !(C)))) */ ;
    defparam i7448_2_lut_3_lut_4_lut.init = 16'h1ef0;
    LUT4 i7462_2_lut_3_lut_4_lut (.A(\pitch_pwm_pulse_length_us[6] ), .B(n52284), 
         .C(\pitch_pwm_pulse_length_us[8] ), .D(\pitch_pwm_pulse_length_us[7] ), 
         .Z(value_out_7__N_154[8])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;
    defparam i7462_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 i24050_3_lut_3_lut (.A(\latched_roll[0] ), .B(\latched_roll[1] ), 
         .C(\latched_roll[3] ), .Z(n34690)) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/angle_controller.v(84[74:86])
    defparam i24050_3_lut_3_lut.init = 16'h6a6a;
    LUT4 i7469_3_lut_4_lut (.A(\pitch_pwm_pulse_length_us[7] ), .B(n52236), 
         .C(\pitch_pwm_pulse_length_us[8] ), .D(\pitch_pwm_pulse_length_us[9] ), 
         .Z(value_out_7__N_154[9])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;
    defparam i7469_3_lut_4_lut.init = 16'h7f80;
    
endmodule
//
// Verilog Description of module \i2c_device_driver(INIT_INTERVAL=16'b01111101000,POLL_INTERVAL=16'b010100) 
//

module \i2c_device_driver(INIT_INTERVAL=16'b01111101000,POLL_INTERVAL=16'b010100)  (sys_clk_N_413, 
            sys_clk, \next_i2c_state_4__N_1055[1] , \next_i2c_device_driver_state[3] , 
            \next_i2c_device_driver_state[2] , \next_i2c_device_driver_state[0] , 
            \next_i2c_device_driver_state[4] , cal_reg_addr, resetn, next_VL53L1X_firm_rdy, 
            \next_i2c_device_driver_return_state[0] , n53885, next_imu_good, 
            \next_i2c_device_driver_return_state[2] , next_VL53L1X_range_mm, 
            next_data_tx_7__N_1032, \next_VL53L1X_data_rdy[7] , next_VL53L1X_chip_id, 
            \next_VL53L1X_data_rdy[6] , \i2c_top_debug[1] , wd_event_active, 
            n52306, \next_VL53L1X_data_rdy[5] , \next_VL53L1X_data_rdy[4] , 
            \next_VL53L1X_data_rdy[3] , \next_VL53L1X_data_rdy[2] , \next_VL53L1X_data_rdy[1] , 
            GND_net, \next_i2c_device_driver_return_state[4] , \next_i2c_device_driver_return_state[3] , 
            \next_i2c_device_driver_return_state[1] , n52205, n52318, 
            \i2c_top_debug[3] , \i2c_top_debug[4] , \next_i2c_device_driver_state[1] , 
            throttle_controller_active, next_imu_data_valid, \next_data_tx_7__N_1032[1] , 
            \i2c_top_debug[0] , \i2c_top_debug[5] , resetn_derived_2, 
            byte_rd_left_5__N_1255, n52142, n27391, n48722, n48829, 
            n52140, i2c2_sdaoen, i2c2_sdao, i2c2_scloen, i2c2_sclo, 
            i2c2_sdai, i2c2_scli, i2c1_sdaoen, i2c1_sdao, i2c1_scloen, 
            i2c1_sclo, i2c1_sdai, i2c1_scli, VCC_net) /* synthesis syn_module_defined=1 */ ;
    input sys_clk_N_413;
    input sys_clk;
    output \next_i2c_state_4__N_1055[1] ;
    output \next_i2c_device_driver_state[3] ;
    output \next_i2c_device_driver_state[2] ;
    output \next_i2c_device_driver_state[0] ;
    output \next_i2c_device_driver_state[4] ;
    output [7:0]cal_reg_addr;
    input resetn;
    output [7:0]next_VL53L1X_firm_rdy;
    output \next_i2c_device_driver_return_state[0] ;
    input n53885;
    output next_imu_good;
    output \next_i2c_device_driver_return_state[2] ;
    output [15:0]next_VL53L1X_range_mm;
    input [7:0]next_data_tx_7__N_1032;
    output \next_VL53L1X_data_rdy[7] ;
    output [15:0]next_VL53L1X_chip_id;
    output \next_VL53L1X_data_rdy[6] ;
    output \i2c_top_debug[1] ;
    output wd_event_active;
    output n52306;
    output \next_VL53L1X_data_rdy[5] ;
    output \next_VL53L1X_data_rdy[4] ;
    output \next_VL53L1X_data_rdy[3] ;
    output \next_VL53L1X_data_rdy[2] ;
    output \next_VL53L1X_data_rdy[1] ;
    input GND_net;
    output \next_i2c_device_driver_return_state[4] ;
    output \next_i2c_device_driver_return_state[3] ;
    output \next_i2c_device_driver_return_state[1] ;
    input n52205;
    input n52318;
    output \i2c_top_debug[3] ;
    output \i2c_top_debug[4] ;
    output \next_i2c_device_driver_state[1] ;
    input throttle_controller_active;
    output next_imu_data_valid;
    input \next_data_tx_7__N_1032[1] ;
    output \i2c_top_debug[0] ;
    output \i2c_top_debug[5] ;
    input resetn_derived_2;
    input byte_rd_left_5__N_1255;
    output n52142;
    input n27391;
    output n48722;
    output n48829;
    input n52140;
    output i2c2_sdaoen;
    output i2c2_sdao;
    output i2c2_scloen;
    output i2c2_sclo;
    input i2c2_sdai;
    input i2c2_scli;
    output i2c1_sdaoen;
    output i2c1_sdao;
    output i2c1_scloen;
    output i2c1_sclo;
    input i2c1_sdai;
    input i2c1_scli;
    input VCC_net;
    
    wire sys_clk_N_413 /* synthesis is_inv_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(82[16:24])
    wire sys_clk /* synthesis SET_AS_NETWORK=sys_clk, is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(220[10:17])
    wire next_addr_7__N_1168 /* synthesis is_clock=1, SET_AS_NETWORK=\I2C_Devices/i2c/next_addr_7__N_1168 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(45[15:24])
    wire i2c2_scli /* synthesis is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_efb_wb.v(34[10:19])
    wire i2c1_scli /* synthesis is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_efb_wb.v(40[10:19])
    wire [16:0]count_sys_clk_for_ms;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(111[15:35])
    wire [16:0]count_sys_clk_for_ms_16__N_857;
    wire [4:0]next_i2c_state_4__N_1090;
    wire [8:0]n7654;
    wire [20:0]master_trigger_count_ms;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(110[15:38])
    
    wire sys_clk_enable_224, n52182;
    wire [20:0]n611;
    wire [7:0]\VL53L1X_data_rx_reg[3] ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(92[15:34])
    
    wire sys_clk_enable_9, n52448;
    wire [7:0]data_rx;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(77[15:22])
    wire [7:0]\VL53L1X_data_rx_reg[2] ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(92[15:34])
    
    wire sys_clk_enable_17, sys_clk_enable_123, n48658, n29, n49469, 
        n52513, n52514, n52515;
    wire [16:0]count_sys_clk_for_ms_16__N_874;
    
    wire n47071, n29_adj_5259, n49454, n53892, n7, n109, n24343, 
        n29_adj_5260, n49457;
    wire [15:0]data_reg;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(73[16:24])
    
    wire n4, resetn_VL53L1X_buffer, n52337, VL53L1X_data_rx_reg_1__4__N_702;
    wire [7:0]data_tx;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(75[15:22])
    
    wire n29_adj_5261, valid_strobe_enable, n46979;
    wire [15:0]VL53L1X_osc_cal_val;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(93[16:35])
    wire [7:0]\VL53L1X_data_rx_reg[5] ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(92[15:34])
    
    wire n30332, VL53L1X_data_rx_reg_7__7__N_473, VL53L1X_data_rx_reg_7__7__N_476, 
        n53891;
    wire [4:0]next_i2c_state_4__N_386;
    wire [4:0]next_return_state_4__N_391;
    wire [31:0]VL53L1X_measurement_period;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(94[16:42])
    
    wire sys_clk_enable_108;
    wire [22:0]next_VL53L1X_measurement_period_31__N_1103;
    
    wire read_write_in;
    wire [8:0]n2485;
    
    wire is_2_byte_reg, sys_clk_enable_73, n15, n52420, n21, n52199;
    wire [15:0]next_data_reg_15__N_362;
    
    wire n8, n14;
    wire [15:0]count_ms;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(82[16:24])
    
    wire n52172, n43843, n8_adj_5262, n49721, n8_adj_5263, n49728, 
        n30336, VL53L1X_data_rx_reg_7__6__N_480, VL53L1X_data_rx_reg_7__6__N_482, 
        n30340, VL53L1X_data_rx_reg_7__5__N_486, VL53L1X_data_rx_reg_7__5__N_488, 
        n46603, n30344, VL53L1X_data_rx_reg_7__4__N_492, VL53L1X_data_rx_reg_7__4__N_494, 
        n30348, VL53L1X_data_rx_reg_7__3__N_498, VL53L1X_data_rx_reg_7__3__N_500, 
        n49722, n30352, VL53L1X_data_rx_reg_7__2__N_504, VL53L1X_data_rx_reg_7__2__N_506, 
        n22, n30356, VL53L1X_data_rx_reg_7__1__N_510, VL53L1X_data_rx_reg_7__1__N_512, 
        n30360, VL53L1X_data_rx_reg_7__0__N_516, VL53L1X_data_rx_reg_7__0__N_518, 
        n30364, VL53L1X_data_rx_reg_6__7__N_522, VL53L1X_data_rx_reg_6__7__N_524, 
        n30368, VL53L1X_data_rx_reg_6__6__N_528, VL53L1X_data_rx_reg_6__6__N_530, 
        n30372, VL53L1X_data_rx_reg_6__5__N_534, VL53L1X_data_rx_reg_6__5__N_536, 
        n52121, n30376, VL53L1X_data_rx_reg_6__4__N_540, VL53L1X_data_rx_reg_6__4__N_542, 
        n52085, n30380, VL53L1X_data_rx_reg_6__3__N_546, VL53L1X_data_rx_reg_6__3__N_548, 
        n52282, n47057, n52136, n30384, VL53L1X_data_rx_reg_6__2__N_552, 
        VL53L1X_data_rx_reg_6__2__N_554, n30388, VL53L1X_data_rx_reg_6__1__N_558, 
        VL53L1X_data_rx_reg_6__1__N_560, n25615;
    wire [2:0]measurement_period_tx_index;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(96[15:42])
    
    wire n51507, n30392, VL53L1X_data_rx_reg_6__0__N_564, VL53L1X_data_rx_reg_6__0__N_566, 
        n51508, n37158, n19, n52137, n30396, VL53L1X_data_rx_reg_5__7__N_570, 
        VL53L1X_data_rx_reg_5__7__N_572, n30400, VL53L1X_data_rx_reg_5__6__N_576, 
        VL53L1X_data_rx_reg_5__6__N_578, n30404, VL53L1X_data_rx_reg_5__5__N_582, 
        VL53L1X_data_rx_reg_5__5__N_584, n30408, VL53L1X_data_rx_reg_5__4__N_588, 
        VL53L1X_data_rx_reg_5__4__N_590, n30412, VL53L1X_data_rx_reg_5__3__N_594, 
        VL53L1X_data_rx_reg_5__3__N_596, n30416, VL53L1X_data_rx_reg_5__2__N_600, 
        VL53L1X_data_rx_reg_5__2__N_602, n30420, VL53L1X_data_rx_reg_5__1__N_606, 
        VL53L1X_data_rx_reg_5__1__N_608, n49495, n30424, VL53L1X_data_rx_reg_5__0__N_612, 
        VL53L1X_data_rx_reg_5__0__N_614, n52484, n30428, VL53L1X_data_rx_reg_4__7__N_618, 
        VL53L1X_data_rx_reg_4__7__N_620, n49720, n30432, VL53L1X_data_rx_reg_4__6__N_624, 
        VL53L1X_data_rx_reg_4__6__N_626, n7_adj_5264, n30436, VL53L1X_data_rx_reg_4__5__N_630, 
        VL53L1X_data_rx_reg_4__5__N_632, n51506, n30440, VL53L1X_data_rx_reg_4__4__N_636, 
        VL53L1X_data_rx_reg_4__4__N_638, n30444, VL53L1X_data_rx_reg_4__3__N_642, 
        VL53L1X_data_rx_reg_4__3__N_644, n30448, VL53L1X_data_rx_reg_4__2__N_648, 
        VL53L1X_data_rx_reg_4__2__N_650, n30452, VL53L1X_data_rx_reg_4__1__N_654, 
        VL53L1X_data_rx_reg_4__1__N_656, n30456, VL53L1X_data_rx_reg_4__0__N_660, 
        VL53L1X_data_rx_reg_4__0__N_662, n30460, VL53L1X_data_rx_reg_1__7__N_682, 
        VL53L1X_data_rx_reg_1__7__N_684;
    wire [15:0]count_ms_15__N_910;
    wire [15:0]count_ms_15__N_894;
    wire [15:0]count_ms_15__N_396;
    
    wire n30464, VL53L1X_data_rx_reg_1__6__N_688, VL53L1X_data_rx_reg_1__6__N_690, 
        n49727, n30468, VL53L1X_data_rx_reg_1__5__N_694, VL53L1X_data_rx_reg_1__5__N_696, 
        n7_adj_5265, n30472, VL53L1X_data_rx_reg_1__4__N_700, n30476, 
        VL53L1X_data_rx_reg_1__3__N_706, VL53L1X_data_rx_reg_1__3__N_708, 
        n30480, VL53L1X_data_rx_reg_1__2__N_712, VL53L1X_data_rx_reg_1__2__N_714, 
        n30484, VL53L1X_data_rx_reg_1__1__N_718, VL53L1X_data_rx_reg_1__1__N_720, 
        n30488, VL53L1X_data_rx_reg_1__0__N_724, VL53L1X_data_rx_reg_1__0__N_726, 
        n30492, VL53L1X_data_rx_reg_0__7__N_730, VL53L1X_data_rx_reg_0__7__N_732, 
        n30496, VL53L1X_data_rx_reg_0__6__N_736, VL53L1X_data_rx_reg_0__6__N_738, 
        n30500, VL53L1X_data_rx_reg_0__5__N_742, VL53L1X_data_rx_reg_0__5__N_744, 
        n30504, VL53L1X_data_rx_reg_0__4__N_748, VL53L1X_data_rx_reg_0__4__N_750, 
        n30508, VL53L1X_data_rx_reg_0__3__N_754, VL53L1X_data_rx_reg_0__3__N_756, 
        n30512, VL53L1X_data_rx_reg_0__2__N_760, VL53L1X_data_rx_reg_0__2__N_762, 
        n30516, VL53L1X_data_rx_reg_0__1__N_766, VL53L1X_data_rx_reg_0__1__N_768, 
        n30520, VL53L1X_data_rx_reg_0__0__N_772, VL53L1X_data_rx_reg_0__0__N_774, 
        n52152, n29_adj_5266, n53873, n7_adj_5267;
    wire [5:0]target_read_count;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(85[15:32])
    
    wire n50875, n52138, n49724, n52526, n52525, n49723, n49725, 
        n52374, n49731, n49729, n49730, n49732, n30613, VL53L1X_data_rx_reg_index_5__N_439, 
        VL53L1X_data_rx_reg_index_5__N_457, n49497, n28220, n19_adj_5268, 
        n20, n21_adj_5269, n52483, n9, n47107, n30, n49468, n30406, 
        n30405, n52360, n30617, VL53L1X_data_rx_reg_index_5__N_442, 
        VL53L1X_data_rx_reg_index_5__N_460, n52351, n52350, n52348, 
        n52347, n52346, n52345, n10, n13, n14_adj_5270, n52344;
    wire [15:0]n44;
    
    wire n52343, n52364, n52363, n52358, n52357, n7_adj_5271, n7250, 
        n52210, n52354, n52352, n76, n52246, n6972, n52574, n52573, 
        n52577, n52576, n52580, n52579, n52583, n52582, n47981, 
        n34032, n14_adj_5272, n47983, n15_adj_5273, n52592, n52591, 
        n52372, n52371, n52370, n47982, n52369, n52368, n52367, 
        n52333, n52366, n52365;
    wire [7:0]\VL53L1X_data_rx_reg[7] ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(92[15:34])
    
    wire n52386, n52384, n15_adj_5274, n52381, n52380, n52377, n52376, 
        n15_adj_5275, n47980, n34018, n27301, n10_adj_5276;
    wire [2:0]next_measurement_period_tx_index;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(97[15:47])
    
    wire n14_adj_5277, n49414, n24, n52440;
    wire [4:0]next_i2c_state_4__N_1050;
    
    wire n37, n53879, n52403, n27913, n52227, n28, n21563, n53;
    wire [5:0]VL53L1X_data_rx_reg_index;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(87[15:40])
    wire [5:0]n6915;
    
    wire n52336, n6974, n48780, VL53L1X_data_rx_reg_index_5__N_463, 
        n6, n52296, n49365, n49547, n43791, n14126, n43792, n52487, 
        n51720, n51721, n49665, n33840, n51722, n7246, n51725, 
        n7_adj_5278, n52314, VL53L1X_data_rx_reg_index_5__N_445, n28_adj_5279, 
        n22284, n52509, n15_adj_5280, n52248, n48104, n29262, n52486, 
        n47394, n50952, n30354, n30353, n52212, sys_clk_enable_242, 
        n53876, n52449, sys_clk_enable_255, n50950, n50951, n52503, 
        n52506, n126, n52154, n19_adj_5281, n28_adj_5282;
    wire [21:0]n2;
    
    wire n30615, n30614, n24_adj_5283, n19_adj_5284, n28_adj_5285, 
        n51817;
    wire [5:0]next_target_read_count_5__N_414;
    
    wire n52274, n125, n52303, n7244;
    wire [6:0]n13173;
    
    wire n51006, n33834, n49511, n52270, n69, n3, n28226, resetn_imu_N_1182, 
        n10_adj_5286, n13_adj_5287, n14_adj_5288, n43790, n52507, 
        n52508, n52412, n52446, n38, n53877, n52444, n52447, one_byte_ready;
    wire [5:0]n23;
    
    wire n28247, n49450, n52203;
    wire [6:0]n13181;
    
    wire n49453, n49456;
    wire [5:0]n13144;
    
    wire n7_adj_5290, n15_adj_5291, n52269, n43789, n52335, n51197, 
        n51199, n52292, n52256;
    wire [63:0]VL53L1X_data_rx_reg_7__7__N_472;
    
    wire n66, n53051, n51131, n51133, n52153, n37517, n51024, 
        n53052, n52460, n51724, n20052, n28_adj_5292, n23389, n51101, 
        n51103, n72, n53050, n52077, n52076, n49226, n52087, n52122, 
        n43788, n7_adj_5293, n7_adj_5294, n14_adj_5295, n14_adj_5296, 
        n47344, n52504, n52505, n52123, n52124, n30346, n30345, 
        n53878, n30350, n30349, n52445;
    wire [7:0]next_data_tx_7__N_1024;
    
    wire n30426, n30425, n30342, n30341, n30338, n30337, n16, 
        n20_adj_5297, n30522, n30521, n52320, n49571, n30518, n30517, 
        n52321, n30334, n30333, n30514, n30513, n52322, n29_adj_5298, 
        n49415, n51099, n51100, n43787, n30510, n30509, n52324;
    wire [20:0]master_trigger_count_ms_20__N_997;
    
    wire n52501, n52502, n14054, n53886, n47760, n52425, n51003, 
        n48098;
    wire [7:0]next_data_tx_7__N_378;
    
    wire n53055, n53054, n53056, n21_adj_5299, n51819, n52231, n43783;
    wire [7:0]next_cal_reg_addr_7__N_1124;
    
    wire n43784, n52271, n49637, n52233, n29_adj_5300, n52218, n52409, 
        n52498, n52499, n7_adj_5301, n7234, n51130, n49625, n49569, 
        n53053, n51129, n52410, n52485, n21_adj_5302, n49478, n52450, 
        n51196, n51195, n22_adj_5303, n49677, n36072, n43986, n1, 
        n52334, n48496, n52177, n3_adj_5304, n23405, n53888, n49535, 
        n52219, n30506, n30505, n52329, n43985, n43984, n43983, 
        n49693, n43982, n30502, n30501, n52330, n30498, n30497, 
        n52331, sys_clk_enable_256, sys_clk_N_413_enable_8, n43981, 
        n30494, n30493, n52332, n30490, n30489, n52042, n18_adj_5312, 
        n6_adj_5313, n30486, n30485, n43786, n43785, n52338, n14_adj_5314, 
        n30482, n30481, n30478, n30477, n43980, n43979, n52078, 
        n19_adj_5319, n52134, n30474, n30473, n52339, n30470, n30469, 
        n46521, n30466, n30465, n28179, n127, n52421, n30_adj_5320, 
        n52283, n52340, n21_adj_5321, n24_adj_5322, n43976;
    wire [22:0]n25;
    
    wire n8_adj_5323, n1_adj_5324, n7_adj_5325, n30462, n30461;
    wire [7:0]next_data_tx_7__N_1032_c;
    
    wire n8_adj_5326, n52040, n52188, n28_adj_5327, n22_adj_5328, 
        n43975, n17827, n43974;
    wire [18:0]n17807;
    
    wire n7240, n43973, n48822, n53890, n43972, n43971, n30458, 
        n30457, n49433, n11_adj_5331, n52209, n22527, n5_adj_5332, 
        n6_adj_5333, n30454, n30453, n48986, n30450, n30449, n43970, 
        n43969, n43968, n43967, n30446, n30445, n30442, n30441, 
        n30438, n30437, n52593, n30434, n30433, n30430, n30429, 
        n30422, n30421, n43966, n43965, n34, n43964, n43963, n43962, 
        n52290, n43961, n43960, n43851, n43959, n52086, n30677, 
        n21625, n49510, n49512, n43956, n43850, n30418, n30417, 
        n52041, n43955, n43954, n43953, n43849, n50826, n30414, 
        n30413, n14_adj_5335, n52135, n52157, n30410, n30409, n49477, 
        n43952, n27, sys_clk_enable_254, n43951, n43848, n43950;
    wire [5:0]next_target_read_count;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(86[15:37])
    
    wire n49101, n43949, n43847, valid_strobe_N_1132, n43846, n43845, 
        n49507, n49508, n51005, n51007, n43805, n43804, n43803, 
        n30402, n30401, n50953, n127_adj_5337, n30398, n30397, n43802, 
        n1_adj_5338, n30394, n30393, rx_from_VL53L1X, n36, n27_adj_5339;
    wire [7:0]i2c_top_debug;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(53[22:35])
    
    wire n45689, n51818, n52201, n33854, n43801, n14_adj_5340, n30390, 
        n30389, n43800, n30386, n30385, n43799, n30619, n30618, 
        n30382, n30381, n30330, n30329, n30328;
    wire [5:0]next_VL53L1X_data_rx_reg_index;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(88[15:45])
    
    wire n30378, n30377, n30374, n30373, n50877, n17_adj_5342, n46519, 
        n48249, n30370, n30369, n30366, n30365, n50878, n43798, 
        n51719, n49472, n48756, n48394, n33, n43797, n30362, n30361, 
        n50879, n50876, n43796, n43794, n43793, n30358, n30357, 
        delay_timer_at_init, go;
    
    FD1S3AY count_sys_clk_for_ms_i0 (.D(count_sys_clk_for_ms_16__N_857[0]), 
            .CK(sys_clk_N_413), .Q(count_sys_clk_for_ms[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam count_sys_clk_for_ms_i0.GSR = "ENABLED";
    FD1S3AX delay_timer_started_488 (.D(n7654[7]), .CK(sys_clk_N_413), .Q(next_i2c_state_4__N_1090[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam delay_timer_started_488.GSR = "ENABLED";
    FD1P3IX master_trigger_count_ms_i0 (.D(n611[0]), .SP(sys_clk_enable_224), 
            .CD(n52182), .CK(sys_clk), .Q(master_trigger_count_ms[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(268[14] 281[12])
    defparam master_trigger_count_ms_i0.GSR = "ENABLED";
    FD1P3DX \VL53L1X_data_rx_reg_3[[7__639  (.D(data_rx[7]), .SP(sys_clk_enable_9), 
            .CK(sys_clk), .CD(n52448), .Q(\VL53L1X_data_rx_reg[3] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_3[[7__639 .GSR = "DISABLED";
    FD1P3DX \VL53L1X_data_rx_reg_3[[6__640  (.D(data_rx[6]), .SP(sys_clk_enable_9), 
            .CK(sys_clk), .CD(n52448), .Q(\VL53L1X_data_rx_reg[3] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_3[[6__640 .GSR = "DISABLED";
    FD1P3DX \VL53L1X_data_rx_reg_3[[5__641  (.D(data_rx[5]), .SP(sys_clk_enable_9), 
            .CK(sys_clk), .CD(n52448), .Q(\VL53L1X_data_rx_reg[3] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_3[[5__641 .GSR = "DISABLED";
    FD1P3DX \VL53L1X_data_rx_reg_3[[4__642  (.D(data_rx[4]), .SP(sys_clk_enable_9), 
            .CK(sys_clk), .CD(n52448), .Q(\VL53L1X_data_rx_reg[3] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_3[[4__642 .GSR = "DISABLED";
    FD1P3DX \VL53L1X_data_rx_reg_3[[3__643  (.D(data_rx[3]), .SP(sys_clk_enable_9), 
            .CK(sys_clk), .CD(n52448), .Q(\VL53L1X_data_rx_reg[3] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_3[[3__643 .GSR = "DISABLED";
    FD1P3DX \VL53L1X_data_rx_reg_3[[2__644  (.D(data_rx[2]), .SP(sys_clk_enable_9), 
            .CK(sys_clk), .CD(n52448), .Q(\VL53L1X_data_rx_reg[3] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_3[[2__644 .GSR = "DISABLED";
    FD1P3DX \VL53L1X_data_rx_reg_3[[1__645  (.D(data_rx[1]), .SP(sys_clk_enable_9), 
            .CK(sys_clk), .CD(n52448), .Q(\VL53L1X_data_rx_reg[3] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_3[[1__645 .GSR = "DISABLED";
    FD1P3DX \VL53L1X_data_rx_reg_3[[0__646  (.D(data_rx[0]), .SP(sys_clk_enable_9), 
            .CK(sys_clk), .CD(n52448), .Q(\VL53L1X_data_rx_reg[3] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_3[[0__646 .GSR = "DISABLED";
    FD1P3DX \VL53L1X_data_rx_reg_2[[7__647  (.D(data_rx[7]), .SP(sys_clk_enable_17), 
            .CK(sys_clk), .CD(n52448), .Q(\VL53L1X_data_rx_reg[2] [7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_2[[7__647 .GSR = "DISABLED";
    FD1P3DX \VL53L1X_data_rx_reg_2[[6__648  (.D(data_rx[6]), .SP(sys_clk_enable_17), 
            .CK(sys_clk), .CD(n52448), .Q(\VL53L1X_data_rx_reg[2] [6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_2[[6__648 .GSR = "DISABLED";
    FD1P3DX \VL53L1X_data_rx_reg_2[[5__649  (.D(data_rx[5]), .SP(sys_clk_enable_17), 
            .CK(sys_clk), .CD(n52448), .Q(\VL53L1X_data_rx_reg[2] [5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_2[[5__649 .GSR = "DISABLED";
    FD1P3DX \VL53L1X_data_rx_reg_2[[4__650  (.D(data_rx[4]), .SP(sys_clk_enable_17), 
            .CK(sys_clk), .CD(n52448), .Q(\VL53L1X_data_rx_reg[2] [4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_2[[4__650 .GSR = "DISABLED";
    FD1P3DX \VL53L1X_data_rx_reg_2[[3__651  (.D(data_rx[3]), .SP(sys_clk_enable_17), 
            .CK(sys_clk), .CD(n52448), .Q(\VL53L1X_data_rx_reg[2] [3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_2[[3__651 .GSR = "DISABLED";
    FD1P3DX \VL53L1X_data_rx_reg_2[[2__652  (.D(data_rx[2]), .SP(sys_clk_enable_17), 
            .CK(sys_clk), .CD(n52448), .Q(\VL53L1X_data_rx_reg[2] [2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_2[[2__652 .GSR = "DISABLED";
    FD1P3DX \VL53L1X_data_rx_reg_2[[1__653  (.D(data_rx[1]), .SP(sys_clk_enable_17), 
            .CK(sys_clk), .CD(n52448), .Q(\VL53L1X_data_rx_reg[2] [1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_2[[1__653 .GSR = "DISABLED";
    FD1P3DX \VL53L1X_data_rx_reg_2[[0__654  (.D(data_rx[0]), .SP(sys_clk_enable_17), 
            .CK(sys_clk), .CD(n52448), .Q(\VL53L1X_data_rx_reg[2] [0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_2[[0__654 .GSR = "DISABLED";
    FD1P3AX VL53L1X_data_rdy__i1 (.D(\VL53L1X_data_rx_reg[3] [0]), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(\next_i2c_state_4__N_1055[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_data_rdy__i1.GSR = "ENABLED";
    PFUMX i38674 (.BLUT(n48658), .ALUT(n29), .C0(\next_i2c_device_driver_state[3] ), 
          .Z(n49469));
    PFUMX i40936 (.BLUT(n52513), .ALUT(n52514), .C0(\next_i2c_device_driver_state[2] ), 
          .Z(n52515));
    LUT4 i25590_2_lut (.A(count_sys_clk_for_ms_16__N_874[0]), .B(n7654[7]), 
         .Z(count_sys_clk_for_ms_16__N_857[0])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(194[14] 219[12])
    defparam i25590_2_lut.init = 16'h8888;
    PFUMX i38659 (.BLUT(n47071), .ALUT(n29_adj_5259), .C0(\next_i2c_device_driver_state[3] ), 
          .Z(n49454));
    LUT4 i23445_4_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), .B(n53892), 
         .C(\next_i2c_device_driver_state[3] ), .D(\next_i2c_device_driver_state[4] ), 
         .Z(n7)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A (B+(C+!(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i23445_4_lut_4_lut.init = 16'h0180;
    LUT4 i25967_4_lut_4_lut (.A(cal_reg_addr[0]), .B(cal_reg_addr[1]), .C(cal_reg_addr[3]), 
         .D(cal_reg_addr[2]), .Z(n109)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A ((C+(D))+!B))) */ ;
    defparam i25967_4_lut_4_lut.init = 16'h0204;
    PFUMX i38662 (.BLUT(n24343), .ALUT(n29_adj_5260), .C0(\next_i2c_device_driver_state[3] ), 
          .Z(n49457));
    LUT4 i1_4_lut_4_lut (.A(n53892), .B(\next_i2c_device_driver_state[0] ), 
         .C(data_reg[8]), .D(\next_i2c_device_driver_state[3] ), .Z(n4)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(B (C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam i1_4_lut_4_lut.init = 16'h6040;
    LUT4 i39566_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52337), 
         .Z(VL53L1X_data_rx_reg_1__4__N_702)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39566_3_lut.init = 16'h5757;
    LUT4 led_data_out_4__I_0_859_Mux_0_i29_4_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n53892), .C(data_tx[0]), .D(\next_i2c_device_driver_state[2] ), 
         .Z(n29_adj_5261)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)))+!A !(B (C (D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam led_data_out_4__I_0_859_Mux_0_i29_4_lut_4_lut.init = 16'h6088;
    FD1S3AX valid_strobe_enable_720 (.D(n52182), .CK(sys_clk), .Q(valid_strobe_enable)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(268[14] 281[12])
    defparam valid_strobe_enable_720.GSR = "ENABLED";
    FD1P3AX VL53L1X_firm_rdy_i0_i0 (.D(\VL53L1X_data_rx_reg[2] [0]), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(next_VL53L1X_firm_rdy[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_firm_rdy_i0_i0.GSR = "ENABLED";
    LUT4 i1_4_lut_4_lut_4_lut (.A(\next_i2c_device_driver_state[4] ), .B(\next_i2c_device_driver_state[0] ), 
         .C(\next_i2c_device_driver_return_state[0] ), .D(n53892), .Z(n46979)) /* synthesis lut_function=(A (C)+!A (B (C+(D))+!B (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam i1_4_lut_4_lut_4_lut.init = 16'hf5e0;
    FD1P3AX VL53L1X_osc_cal_val_i0_i0 (.D(\VL53L1X_data_rx_reg[5] [0]), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(VL53L1X_osc_cal_val[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_osc_cal_val_i0_i0.GSR = "ENABLED";
    FD1S1D i19660 (.D(n53885), .CK(VL53L1X_data_rx_reg_7__7__N_473), .CD(VL53L1X_data_rx_reg_7__7__N_476), 
           .Q(n30332));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19660.GSR = "DISABLED";
    FD1S3IX i2c_state__i1 (.D(next_i2c_state_4__N_386[0]), .CK(sys_clk), 
            .CD(n53891), .Q(\next_i2c_device_driver_state[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam i2c_state__i1.GSR = "ENABLED";
    FD1S3IX return_state__i1 (.D(next_return_state_4__N_391[0]), .CK(sys_clk), 
            .CD(n53891), .Q(\next_i2c_device_driver_return_state[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam return_state__i1.GSR = "ENABLED";
    FD1P3IX VL53L1X_measurement_period__i0 (.D(next_VL53L1X_measurement_period_31__N_1103[2]), 
            .SP(sys_clk_enable_108), .CD(n53891), .CK(sys_clk), .Q(VL53L1X_measurement_period[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam VL53L1X_measurement_period__i0.GSR = "ENABLED";
    FD1S3IX read_write_in_729 (.D(n2485[3]), .CK(sys_clk), .CD(n53891), 
            .Q(read_write_in)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam read_write_in_729.GSR = "ENABLED";
    FD1S3IX imu_good_736 (.D(n2485[5]), .CK(sys_clk), .CD(n53891), .Q(next_imu_good)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam imu_good_736.GSR = "ENABLED";
    FD1S3IX is_2_byte_reg_739 (.D(n2485[2]), .CK(sys_clk), .CD(n53891), 
            .Q(is_2_byte_reg)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam is_2_byte_reg_739.GSR = "ENABLED";
    FD1P3JX cal_reg_addr_i0 (.D(n15), .SP(sys_clk_enable_73), .PD(n53891), 
            .CK(sys_clk), .Q(cal_reg_addr[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam cal_reg_addr_i0.GSR = "ENABLED";
    FD1S3AY resetn_VL53L1X_buffer_742 (.D(n7654[4]), .CK(sys_clk), .Q(resetn_VL53L1X_buffer)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam resetn_VL53L1X_buffer_742.GSR = "ENABLED";
    FD1P3IX master_trigger_count_ms_i2 (.D(n611[2]), .SP(sys_clk_enable_224), 
            .CD(n52182), .CK(sys_clk), .Q(master_trigger_count_ms[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(268[14] 281[12])
    defparam master_trigger_count_ms_i2.GSR = "ENABLED";
    LUT4 i39213_3_lut_rep_263_4_lut (.A(n52420), .B(data_tx[6]), .C(\next_i2c_device_driver_state[3] ), 
         .D(n21), .Z(n52199)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam i39213_3_lut_rep_263_4_lut.init = 16'h8f80;
    FD1S3IX data_reg__i0 (.D(next_data_reg_15__N_362[0]), .CK(sys_clk), 
            .CD(n53891), .Q(data_reg[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam data_reg__i0.GSR = "ENABLED";
    LUT4 led_data_out_4__I_0_859_Mux_6_i14_4_lut_4_lut_4_lut (.A(n53892), 
         .B(\next_i2c_device_driver_state[2] ), .C(\next_i2c_device_driver_state[0] ), 
         .D(n8), .Z(n14)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B+!(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam led_data_out_4__I_0_859_Mux_6_i14_4_lut_4_lut_4_lut.init = 16'h1908;
    FD1P3IX count_ms_i0 (.D(n43843), .SP(count_sys_clk_for_ms[16]), .CD(n52172), 
            .CK(sys_clk_N_413), .Q(count_ms[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam count_ms_i0.GSR = "ENABLED";
    LUT4 i38926_4_lut_4_lut_4_lut (.A(n53892), .B(\next_i2c_device_driver_state[2] ), 
         .C(\next_i2c_device_driver_state[0] ), .D(n8_adj_5262), .Z(n49721)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B+!(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i38926_4_lut_4_lut_4_lut.init = 16'h1908;
    LUT4 i38933_4_lut_4_lut_4_lut (.A(n53892), .B(\next_i2c_device_driver_state[2] ), 
         .C(\next_i2c_device_driver_state[0] ), .D(n8_adj_5263), .Z(n49728)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B+!(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i38933_4_lut_4_lut_4_lut.init = 16'h1908;
    FD1S1D i19664 (.D(n53885), .CK(VL53L1X_data_rx_reg_7__6__N_480), .CD(VL53L1X_data_rx_reg_7__6__N_482), 
           .Q(n30336));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19664.GSR = "DISABLED";
    FD1S1D i19668 (.D(n53885), .CK(VL53L1X_data_rx_reg_7__5__N_486), .CD(VL53L1X_data_rx_reg_7__5__N_488), 
           .Q(n30340));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19668.GSR = "DISABLED";
    LUT4 i21_4_lut_4_lut_4_lut (.A(n53892), .B(\next_i2c_device_driver_state[0] ), 
         .C(\next_i2c_device_driver_return_state[0] ), .D(\next_i2c_device_driver_state[4] ), 
         .Z(n46603)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C+(D))+!B !(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i21_4_lut_4_lut_4_lut.init = 16'h6651;
    FD1S1D i19672 (.D(n53885), .CK(VL53L1X_data_rx_reg_7__4__N_492), .CD(VL53L1X_data_rx_reg_7__4__N_494), 
           .Q(n30344));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19672.GSR = "DISABLED";
    FD1S1D i19676 (.D(n53885), .CK(VL53L1X_data_rx_reg_7__3__N_498), .CD(VL53L1X_data_rx_reg_7__3__N_500), 
           .Q(n30348));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19676.GSR = "DISABLED";
    LUT4 i38927_3_lut_3_lut_4_lut (.A(n53892), .B(\next_i2c_device_driver_state[2] ), 
         .C(\next_i2c_device_driver_state[0] ), .D(data_reg[7]), .Z(n49722)) /* synthesis lut_function=(A (B (C))+!A (((D)+!C)+!B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i38927_3_lut_3_lut_4_lut.init = 16'hd595;
    FD1S1D i19680 (.D(n53885), .CK(VL53L1X_data_rx_reg_7__2__N_504), .CD(VL53L1X_data_rx_reg_7__2__N_506), 
           .Q(n30352));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19680.GSR = "DISABLED";
    LUT4 i26743_4_lut_4_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n53892), .C(\next_i2c_device_driver_state[2] ), .D(data_reg[5]), 
         .Z(n22)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(B (C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam i26743_4_lut_4_lut_4_lut.init = 16'h6040;
    FD1S1D i19684 (.D(n53885), .CK(VL53L1X_data_rx_reg_7__1__N_510), .CD(VL53L1X_data_rx_reg_7__1__N_512), 
           .Q(n30356));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19684.GSR = "DISABLED";
    FD1S1D i19688 (.D(n53885), .CK(VL53L1X_data_rx_reg_7__0__N_516), .CD(VL53L1X_data_rx_reg_7__0__N_518), 
           .Q(n30360));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19688.GSR = "DISABLED";
    FD1S1D i19692 (.D(n53885), .CK(VL53L1X_data_rx_reg_6__7__N_522), .CD(VL53L1X_data_rx_reg_6__7__N_524), 
           .Q(n30364));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19692.GSR = "DISABLED";
    FD1S1D i19696 (.D(n53885), .CK(VL53L1X_data_rx_reg_6__6__N_528), .CD(VL53L1X_data_rx_reg_6__6__N_530), 
           .Q(n30368));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19696.GSR = "DISABLED";
    FD1S1D i19700 (.D(n53885), .CK(VL53L1X_data_rx_reg_6__5__N_534), .CD(VL53L1X_data_rx_reg_6__5__N_536), 
           .Q(n30372));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19700.GSR = "DISABLED";
    LUT4 n7_bdd_3_lut_40892_3_lut_4_lut (.A(\next_i2c_device_driver_state[2] ), 
         .B(\next_i2c_device_driver_state[0] ), .C(\next_i2c_device_driver_state[3] ), 
         .D(n53892), .Z(n52121)) /* synthesis lut_function=(!(A (B (C (D)))+!A !(B+((D)+!C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam n7_bdd_3_lut_40892_3_lut_4_lut.init = 16'h7fef;
    FD1S1D i19704 (.D(n53885), .CK(VL53L1X_data_rx_reg_6__4__N_540), .CD(VL53L1X_data_rx_reg_6__4__N_542), 
           .Q(n30376));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19704.GSR = "DISABLED";
    LUT4 n24200_bdd_4_lut_4_lut (.A(\next_i2c_device_driver_state[2] ), .B(n53892), 
         .C(\next_i2c_device_driver_state[3] ), .D(\next_i2c_device_driver_state[0] ), 
         .Z(n52085)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+((D)+!C))) */ ;
    defparam n24200_bdd_4_lut_4_lut.init = 16'hfdef;
    FD1S1D i19708 (.D(n53885), .CK(VL53L1X_data_rx_reg_6__3__N_546), .CD(VL53L1X_data_rx_reg_6__3__N_548), 
           .Q(n30380));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19708.GSR = "DISABLED";
    LUT4 data_reg_6__bdd_4_lut (.A(data_reg[6]), .B(n52282), .C(n47057), 
         .D(\next_i2c_device_driver_state[3] ), .Z(n52136)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A !((D)+!C)) */ ;
    defparam data_reg_6__bdd_4_lut.init = 16'h88f0;
    FD1S1D i19712 (.D(n53885), .CK(VL53L1X_data_rx_reg_6__2__N_552), .CD(VL53L1X_data_rx_reg_6__2__N_554), 
           .Q(n30384));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19712.GSR = "DISABLED";
    FD1S1D i19716 (.D(n53885), .CK(VL53L1X_data_rx_reg_6__1__N_558), .CD(VL53L1X_data_rx_reg_6__1__N_560), 
           .Q(n30388));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19716.GSR = "DISABLED";
    LUT4 i15152_3_lut_4_lut_4_lut_4_lut (.A(n53892), .B(\next_i2c_device_driver_state[0] ), 
         .C(\next_i2c_device_driver_state[3] ), .D(\next_i2c_device_driver_state[2] ), 
         .Z(n25615)) /* synthesis lut_function=(A (B+(C+(D)))+!A !(B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam i15152_3_lut_4_lut_4_lut_4_lut.init = 16'hbfb8;
    LUT4 measurement_period_tx_index_0__bdd_3_lut_40857 (.A(VL53L1X_measurement_period[2]), 
         .B(measurement_period_tx_index[1]), .C(VL53L1X_measurement_period[18]), 
         .Z(n51507)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam measurement_period_tx_index_0__bdd_3_lut_40857.init = 16'he2e2;
    FD1S1D i19720 (.D(n53885), .CK(VL53L1X_data_rx_reg_6__0__N_564), .CD(VL53L1X_data_rx_reg_6__0__N_566), 
           .Q(n30392));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19720.GSR = "DISABLED";
    LUT4 n51508_bdd_4_lut (.A(n51508), .B(n37158), .C(n19), .D(n53892), 
         .Z(n52137)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A !((D)+!C)) */ ;
    defparam n51508_bdd_4_lut.init = 16'h88f0;
    FD1S1D i19724 (.D(n53885), .CK(VL53L1X_data_rx_reg_5__7__N_570), .CD(VL53L1X_data_rx_reg_5__7__N_572), 
           .Q(n30396));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19724.GSR = "DISABLED";
    FD1S1D i19728 (.D(n53885), .CK(VL53L1X_data_rx_reg_5__6__N_576), .CD(VL53L1X_data_rx_reg_5__6__N_578), 
           .Q(n30400));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19728.GSR = "DISABLED";
    FD1S1D i19732 (.D(n53885), .CK(VL53L1X_data_rx_reg_5__5__N_582), .CD(VL53L1X_data_rx_reg_5__5__N_584), 
           .Q(n30404));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19732.GSR = "DISABLED";
    FD1S1D i19736 (.D(n53885), .CK(VL53L1X_data_rx_reg_5__4__N_588), .CD(VL53L1X_data_rx_reg_5__4__N_590), 
           .Q(n30408));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19736.GSR = "DISABLED";
    FD1S1D i19740 (.D(n53885), .CK(VL53L1X_data_rx_reg_5__3__N_594), .CD(VL53L1X_data_rx_reg_5__3__N_596), 
           .Q(n30412));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19740.GSR = "DISABLED";
    FD1S1D i19744 (.D(n53885), .CK(VL53L1X_data_rx_reg_5__2__N_600), .CD(VL53L1X_data_rx_reg_5__2__N_602), 
           .Q(n30416));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19744.GSR = "DISABLED";
    FD1S1D i19748 (.D(n53885), .CK(VL53L1X_data_rx_reg_5__1__N_606), .CD(VL53L1X_data_rx_reg_5__1__N_608), 
           .Q(n30420));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19748.GSR = "DISABLED";
    LUT4 i38700_4_lut_4_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n53892), .C(\next_i2c_device_driver_state[2] ), .D(\next_i2c_device_driver_return_state[2] ), 
         .Z(n49495)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i38700_4_lut_4_lut_4_lut.init = 16'h1f18;
    FD1S1D i19752 (.D(n53885), .CK(VL53L1X_data_rx_reg_5__0__N_612), .CD(VL53L1X_data_rx_reg_5__0__N_614), 
           .Q(n30424));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19752.GSR = "DISABLED";
    LUT4 led_data_out_4__I_0_862_Mux_1_i22_4_lut_then_4_lut (.A(\next_i2c_device_driver_state[2] ), 
         .B(\next_i2c_device_driver_state[3] ), .C(n53892), .D(\next_i2c_device_driver_state[0] ), 
         .Z(n52484)) /* synthesis lut_function=(A (B+!(C (D)+!C !(D)))+!A !(B ((D)+!C)+!B (C (D)+!C !(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam led_data_out_4__I_0_862_Mux_1_i22_4_lut_then_4_lut.init = 16'h8bf8;
    FD1S1D i19756 (.D(n53885), .CK(VL53L1X_data_rx_reg_4__7__N_618), .CD(VL53L1X_data_rx_reg_4__7__N_620), 
           .Q(n30428));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19756.GSR = "DISABLED";
    LUT4 i38925_4_lut_4_lut_4_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n53892), .C(data_reg[7]), .D(\next_i2c_device_driver_state[2] ), 
         .Z(n49720)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i38925_4_lut_4_lut_4_lut_4_lut.init = 16'h1170;
    FD1S1D i19760 (.D(n53885), .CK(VL53L1X_data_rx_reg_4__6__N_624), .CD(VL53L1X_data_rx_reg_4__6__N_626), 
           .Q(n30432));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19760.GSR = "DISABLED";
    LUT4 led_data_out_4__I_0_858_Mux_6_i7_4_lut_4_lut_4_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n53892), .C(data_reg[6]), .D(\next_i2c_device_driver_state[2] ), 
         .Z(n7_adj_5264)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B ((D)+!C)+!B !(C+(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam led_data_out_4__I_0_858_Mux_6_i7_4_lut_4_lut_4_lut_4_lut.init = 16'h1170;
    FD1S1D i19764 (.D(n53885), .CK(VL53L1X_data_rx_reg_4__5__N_630), .CD(VL53L1X_data_rx_reg_4__5__N_632), 
           .Q(n30436));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19764.GSR = "DISABLED";
    LUT4 measurement_period_tx_index_0__bdd_2_lut_40856 (.A(measurement_period_tx_index[1]), 
         .B(VL53L1X_measurement_period[10]), .Z(n51506)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam measurement_period_tx_index_0__bdd_2_lut_40856.init = 16'h4444;
    FD1S1D i19768 (.D(n53885), .CK(VL53L1X_data_rx_reg_4__4__N_636), .CD(VL53L1X_data_rx_reg_4__4__N_638), 
           .Q(n30440));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19768.GSR = "DISABLED";
    FD1S1D i19772 (.D(n53885), .CK(VL53L1X_data_rx_reg_4__3__N_642), .CD(VL53L1X_data_rx_reg_4__3__N_644), 
           .Q(n30444));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19772.GSR = "DISABLED";
    FD1S1D i19776 (.D(n53885), .CK(VL53L1X_data_rx_reg_4__2__N_648), .CD(VL53L1X_data_rx_reg_4__2__N_650), 
           .Q(n30448));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19776.GSR = "DISABLED";
    FD1S1D i19780 (.D(n53885), .CK(VL53L1X_data_rx_reg_4__1__N_654), .CD(VL53L1X_data_rx_reg_4__1__N_656), 
           .Q(n30452));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19780.GSR = "DISABLED";
    FD1S1D i19784 (.D(n53885), .CK(VL53L1X_data_rx_reg_4__0__N_660), .CD(VL53L1X_data_rx_reg_4__0__N_662), 
           .Q(n30456));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19784.GSR = "DISABLED";
    FD1S1D i19788 (.D(n53885), .CK(VL53L1X_data_rx_reg_1__7__N_682), .CD(VL53L1X_data_rx_reg_1__7__N_684), 
           .Q(n30460));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19788.GSR = "DISABLED";
    LUT4 count_ms_15__I_0_875_i6_3_lut (.A(count_ms_15__N_910[4]), .B(count_ms_15__N_894[5]), 
         .C(n7654[7]), .Z(count_ms_15__N_396[5])) /* synthesis lut_function=(A (B (C))+!A (B+!(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(194[14] 219[12])
    defparam count_ms_15__I_0_875_i6_3_lut.init = 16'hc5c5;
    FD1S1D i19792 (.D(n53885), .CK(VL53L1X_data_rx_reg_1__6__N_688), .CD(VL53L1X_data_rx_reg_1__6__N_690), 
           .Q(n30464));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19792.GSR = "DISABLED";
    LUT4 i38932_4_lut_4_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n53892), .C(\next_i2c_device_driver_state[2] ), .D(data_reg[2]), 
         .Z(n49727)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i38932_4_lut_4_lut_4_lut.init = 16'h1f18;
    FD1S1D i19796 (.D(n53885), .CK(VL53L1X_data_rx_reg_1__5__N_694), .CD(VL53L1X_data_rx_reg_1__5__N_696), 
           .Q(n30468));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19796.GSR = "DISABLED";
    LUT4 led_data_out_4__I_0_858_Mux_5_i7_4_lut_4_lut_4_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n53892), .C(\next_i2c_device_driver_state[2] ), .D(data_reg[5]), 
         .Z(n7_adj_5265)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam led_data_out_4__I_0_858_Mux_5_i7_4_lut_4_lut_4_lut_4_lut.init = 16'h1710;
    FD1S1D i19800 (.D(n53885), .CK(VL53L1X_data_rx_reg_1__4__N_700), .CD(VL53L1X_data_rx_reg_1__4__N_702), 
           .Q(n30472));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19800.GSR = "DISABLED";
    FD1S1D i19804 (.D(n53885), .CK(VL53L1X_data_rx_reg_1__3__N_706), .CD(VL53L1X_data_rx_reg_1__3__N_708), 
           .Q(n30476));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19804.GSR = "DISABLED";
    FD1S1D i19808 (.D(n53885), .CK(VL53L1X_data_rx_reg_1__2__N_712), .CD(VL53L1X_data_rx_reg_1__2__N_714), 
           .Q(n30480));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19808.GSR = "DISABLED";
    FD1S1D i19812 (.D(n53885), .CK(VL53L1X_data_rx_reg_1__1__N_718), .CD(VL53L1X_data_rx_reg_1__1__N_720), 
           .Q(n30484));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19812.GSR = "DISABLED";
    FD1S1D i19816 (.D(n53885), .CK(VL53L1X_data_rx_reg_1__0__N_724), .CD(VL53L1X_data_rx_reg_1__0__N_726), 
           .Q(n30488));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19816.GSR = "DISABLED";
    FD1S1D i19820 (.D(n53885), .CK(VL53L1X_data_rx_reg_0__7__N_730), .CD(VL53L1X_data_rx_reg_0__7__N_732), 
           .Q(n30492));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19820.GSR = "DISABLED";
    FD1S1D i19824 (.D(n53885), .CK(VL53L1X_data_rx_reg_0__6__N_736), .CD(VL53L1X_data_rx_reg_0__6__N_738), 
           .Q(n30496));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19824.GSR = "DISABLED";
    FD1S1D i19828 (.D(n53885), .CK(VL53L1X_data_rx_reg_0__5__N_742), .CD(VL53L1X_data_rx_reg_0__5__N_744), 
           .Q(n30500));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19828.GSR = "DISABLED";
    FD1S1D i19832 (.D(n53885), .CK(VL53L1X_data_rx_reg_0__4__N_748), .CD(VL53L1X_data_rx_reg_0__4__N_750), 
           .Q(n30504));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19832.GSR = "DISABLED";
    FD1S1D i19836 (.D(n53885), .CK(VL53L1X_data_rx_reg_0__3__N_754), .CD(VL53L1X_data_rx_reg_0__3__N_756), 
           .Q(n30508));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19836.GSR = "DISABLED";
    FD1S1D i19840 (.D(n53885), .CK(VL53L1X_data_rx_reg_0__2__N_760), .CD(VL53L1X_data_rx_reg_0__2__N_762), 
           .Q(n30512));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19840.GSR = "DISABLED";
    FD1S1D i19844 (.D(n53885), .CK(VL53L1X_data_rx_reg_0__1__N_766), .CD(VL53L1X_data_rx_reg_0__1__N_768), 
           .Q(n30516));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19844.GSR = "DISABLED";
    FD1S1D i19848 (.D(n53885), .CK(VL53L1X_data_rx_reg_0__0__N_772), .CD(VL53L1X_data_rx_reg_0__0__N_774), 
           .Q(n30520));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19848.GSR = "DISABLED";
    LUT4 n52152_bdd_4_lut (.A(n52152), .B(\next_i2c_device_driver_state[2] ), 
         .C(n29_adj_5266), .D(\next_i2c_device_driver_state[3] ), .Z(n53873)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C (D))) */ ;
    defparam n52152_bdd_4_lut.init = 16'hf088;
    LUT4 led_data_out_4__I_0_860_Mux_2_i7_3_lut_4_lut_4_lut (.A(next_VL53L1X_firm_rdy[0]), 
         .B(\next_i2c_device_driver_state[0] ), .C(n53892), .D(\next_i2c_device_driver_state[2] ), 
         .Z(n7_adj_5267)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A (B ((D)+!C)+!B (C+!(D))))) */ ;
    defparam led_data_out_4__I_0_860_Mux_2_i7_3_lut_4_lut_4_lut.init = 16'h01c0;
    LUT4 n13_bdd_4_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), .B(n53892), 
         .C(target_read_count[1]), .D(\next_i2c_device_driver_state[2] ), 
         .Z(n50875)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam n13_bdd_4_lut_4_lut.init = 16'hf0c4;
    LUT4 next_i2c_device_driver_return_state_2__bdd_4_lut_4_lut (.A(\next_i2c_device_driver_return_state[2] ), 
         .B(n53892), .C(\next_i2c_device_driver_state[0] ), .D(\next_i2c_device_driver_state[2] ), 
         .Z(n52138)) /* synthesis lut_function=(A (B (D)+!B (C))+!A (B (D))) */ ;
    defparam next_i2c_device_driver_return_state_2__bdd_4_lut_4_lut.init = 16'hec20;
    PFUMX i38929 (.BLUT(n49720), .ALUT(n49721), .C0(\next_i2c_device_driver_state[3] ), 
          .Z(n49724));
    LUT4 i1_4_lut_4_lut_then_3_lut (.A(n53892), .B(\next_i2c_device_driver_state[0] ), 
         .C(\next_i2c_device_driver_state[3] ), .Z(n52526)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i1_4_lut_4_lut_then_3_lut.init = 16'h0101;
    LUT4 i1_4_lut_4_lut_else_3_lut (.A(n53892), .B(\next_i2c_device_driver_state[3] ), 
         .C(\next_i2c_device_driver_state[4] ), .Z(n52525)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i1_4_lut_4_lut_else_3_lut.init = 16'h4040;
    PFUMX i38930 (.BLUT(n49722), .ALUT(n49723), .C0(\next_i2c_device_driver_state[3] ), 
          .Z(n49725));
    FD1P3AX VL53L1X_range_mm_i0_i0 (.D(n52374), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(next_VL53L1X_range_mm[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_range_mm_i0_i0.GSR = "ENABLED";
    FD1P3IX master_trigger_count_ms_i1 (.D(n611[1]), .SP(sys_clk_enable_224), 
            .CD(n52182), .CK(sys_clk), .Q(master_trigger_count_ms[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(268[14] 281[12])
    defparam master_trigger_count_ms_i1.GSR = "ENABLED";
    PFUMX i38936 (.BLUT(n49727), .ALUT(n49728), .C0(\next_i2c_device_driver_state[3] ), 
          .Z(n49731));
    PFUMX i38937 (.BLUT(n49729), .ALUT(n49730), .C0(\next_i2c_device_driver_state[3] ), 
          .Z(n49732));
    LUT4 count_ms_15__I_0_875_i5_3_lut (.A(count_ms_15__N_910[4]), .B(count_ms_15__N_894[4]), 
         .C(n7654[7]), .Z(count_ms_15__N_396[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(194[14] 219[12])
    defparam count_ms_15__I_0_875_i5_3_lut.init = 16'hcaca;
    FD1S1D i19941 (.D(n53885), .CK(VL53L1X_data_rx_reg_index_5__N_439), 
           .CD(VL53L1X_data_rx_reg_index_5__N_457), .Q(n30613));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(229[14] 230[75])
    defparam i19941.GSR = "DISABLED";
    LUT4 i39725_2_lut (.A(measurement_period_tx_index[2]), .B(\next_i2c_device_driver_state[0] ), 
         .Z(n37158)) /* synthesis lut_function=(!(A+(B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam i39725_2_lut.init = 16'h1111;
    PFUMX led_data_out_4__I_0_862_Mux_2_i31 (.BLUT(n49497), .ALUT(n28220), 
          .C0(\next_i2c_device_driver_state[4] ), .Z(next_return_state_4__N_391[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;
    PFUMX led_data_out_4__I_0_859_Mux_5_i21 (.BLUT(n19_adj_5268), .ALUT(n20), 
          .C0(n53892), .Z(n21_adj_5269)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;
    LUT4 led_data_out_4__I_0_862_Mux_1_i22_4_lut_else_4_lut (.A(\next_i2c_device_driver_state[2] ), 
         .B(\next_i2c_device_driver_state[3] ), .C(n53892), .D(\next_i2c_device_driver_state[0] ), 
         .Z(n52483)) /* synthesis lut_function=(!(A (B+(C (D)+!C !(D)))+!A (B ((D)+!C)+!B (C (D)+!C !(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam led_data_out_4__I_0_862_Mux_1_i22_4_lut_else_4_lut.init = 16'h0370;
    PFUMX i38673 (.BLUT(n9), .ALUT(n47107), .C0(n30), .Z(n49468));
    LUT4 i19735_3_lut_rep_424 (.A(n30406), .B(n30405), .C(n30404), .Z(n52360)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19735_3_lut_rep_424.init = 16'hcaca;
    FD1S1D i19945 (.D(n53885), .CK(VL53L1X_data_rx_reg_index_5__N_442), 
           .CD(VL53L1X_data_rx_reg_index_5__N_460), .Q(n30617));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(229[14] 230[75])
    defparam i19945.GSR = "DISABLED";
    FD1P3AX VL53L1X_osc_cal_val_i0_i15 (.D(n52351), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(VL53L1X_osc_cal_val[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_osc_cal_val_i0_i15.GSR = "ENABLED";
    FD1P3AX VL53L1X_osc_cal_val_i0_i14 (.D(n52350), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(VL53L1X_osc_cal_val[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_osc_cal_val_i0_i14.GSR = "ENABLED";
    FD1P3AX VL53L1X_osc_cal_val_i0_i13 (.D(n52348), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(VL53L1X_osc_cal_val[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_osc_cal_val_i0_i13.GSR = "ENABLED";
    FD1P3AX VL53L1X_osc_cal_val_i0_i12 (.D(n52347), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(VL53L1X_osc_cal_val[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_osc_cal_val_i0_i12.GSR = "ENABLED";
    FD1P3AX VL53L1X_osc_cal_val_i0_i11 (.D(n52346), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(VL53L1X_osc_cal_val[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_osc_cal_val_i0_i11.GSR = "ENABLED";
    FD1P3AX VL53L1X_osc_cal_val_i0_i10 (.D(n52345), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(VL53L1X_osc_cal_val[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_osc_cal_val_i0_i10.GSR = "ENABLED";
    PFUMX led_data_out_4__I_0_862_Mux_1_i14 (.BLUT(n10), .ALUT(n13), .C0(\next_i2c_device_driver_state[2] ), 
          .Z(n14_adj_5270)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;
    FD1P3AX VL53L1X_osc_cal_val_i0_i9 (.D(n52344), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(VL53L1X_osc_cal_val[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_osc_cal_val_i0_i9.GSR = "ENABLED";
    LUT4 i25970_4_lut (.A(count_ms[3]), .B(n7654[7]), .C(n44[3]), .D(count_sys_clk_for_ms[16]), 
         .Z(count_ms_15__N_396[3])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(194[14] 219[12])
    defparam i25970_4_lut.init = 16'hc088;
    FD1P3AX VL53L1X_osc_cal_val_i0_i8 (.D(n52343), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(VL53L1X_osc_cal_val[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_osc_cal_val_i0_i8.GSR = "ENABLED";
    FD1P3AX VL53L1X_osc_cal_val_i0_i7 (.D(n52364), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(VL53L1X_osc_cal_val[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_osc_cal_val_i0_i7.GSR = "ENABLED";
    FD1P3AX VL53L1X_osc_cal_val_i0_i6 (.D(n52363), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(VL53L1X_osc_cal_val[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_osc_cal_val_i0_i6.GSR = "ENABLED";
    FD1P3AX VL53L1X_osc_cal_val_i0_i5 (.D(n52360), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(VL53L1X_osc_cal_val[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_osc_cal_val_i0_i5.GSR = "ENABLED";
    FD1P3AX VL53L1X_osc_cal_val_i0_i4 (.D(n52358), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(VL53L1X_osc_cal_val[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_osc_cal_val_i0_i4.GSR = "ENABLED";
    FD1P3AX VL53L1X_osc_cal_val_i0_i3 (.D(n52357), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(VL53L1X_osc_cal_val[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_osc_cal_val_i0_i3.GSR = "ENABLED";
    LUT4 i4_4_lut (.A(n7_adj_5271), .B(n7250), .C(\next_i2c_device_driver_state[0] ), 
         .D(n52210), .Z(n7654[6])) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i4_4_lut.init = 16'h8000;
    FD1P3AX VL53L1X_osc_cal_val_i0_i2 (.D(n52354), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(VL53L1X_osc_cal_val[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_osc_cal_val_i0_i2.GSR = "ENABLED";
    FD1P3AX VL53L1X_osc_cal_val_i0_i1 (.D(n52352), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(VL53L1X_osc_cal_val[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_osc_cal_val_i0_i1.GSR = "ENABLED";
    FD1P3AX VL53L1X_firm_rdy_i0_i7 (.D(\VL53L1X_data_rx_reg[2] [7]), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(next_VL53L1X_firm_rdy[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_firm_rdy_i0_i7.GSR = "ENABLED";
    FD1P3AX VL53L1X_firm_rdy_i0_i6 (.D(\VL53L1X_data_rx_reg[2] [6]), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(next_VL53L1X_firm_rdy[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_firm_rdy_i0_i6.GSR = "ENABLED";
    LUT4 n76_bdd_4_lut (.A(n76), .B(n7), .C(\next_i2c_device_driver_state[2] ), 
         .D(n52246), .Z(n6972)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam n76_bdd_4_lut.init = 16'hca00;
    LUT4 n34957_bdd_4_lut_40902_4_lut_then_4_lut (.A(next_data_tx_7__N_1032[3]), 
         .B(\next_i2c_device_driver_state[0] ), .C(n53892), .D(data_tx[3]), 
         .Z(n52574)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C))+!A ((C+!(D))+!B))) */ ;
    defparam n34957_bdd_4_lut_40902_4_lut_then_4_lut.init = 16'h0e02;
    LUT4 n34957_bdd_4_lut_40902_4_lut_else_4_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n53892), .C(data_tx[3]), .Z(n52573)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam n34957_bdd_4_lut_40902_4_lut_else_4_lut.init = 16'h7070;
    LUT4 n34957_bdd_4_lut_40903_4_lut_then_4_lut (.A(next_data_tx_7__N_1032[5]), 
         .B(\next_i2c_device_driver_state[0] ), .C(n53892), .D(data_tx[5]), 
         .Z(n52577)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C))+!A ((C+!(D))+!B))) */ ;
    defparam n34957_bdd_4_lut_40903_4_lut_then_4_lut.init = 16'h0e02;
    LUT4 n34957_bdd_4_lut_40903_4_lut_else_4_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n53892), .C(data_tx[5]), .Z(n52576)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam n34957_bdd_4_lut_40903_4_lut_else_4_lut.init = 16'h7070;
    LUT4 n34957_bdd_4_lut_40901_4_lut_then_4_lut (.A(next_data_tx_7__N_1032[7]), 
         .B(\next_i2c_device_driver_state[0] ), .C(n53892), .D(data_tx[7]), 
         .Z(n52580)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C))+!A ((C+!(D))+!B))) */ ;
    defparam n34957_bdd_4_lut_40901_4_lut_then_4_lut.init = 16'h0e02;
    LUT4 n34957_bdd_4_lut_40901_4_lut_else_4_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n53892), .C(data_tx[7]), .Z(n52579)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam n34957_bdd_4_lut_40901_4_lut_else_4_lut.init = 16'h7070;
    LUT4 n34957_bdd_4_lut_4_lut_then_4_lut (.A(next_data_tx_7__N_1032[2]), 
         .B(\next_i2c_device_driver_state[0] ), .C(n53892), .D(data_tx[2]), 
         .Z(n52583)) /* synthesis lut_function=(!(A (B (C+!(D))+!B (C))+!A ((C+!(D))+!B))) */ ;
    defparam n34957_bdd_4_lut_4_lut_then_4_lut.init = 16'h0e02;
    LUT4 n34957_bdd_4_lut_4_lut_else_4_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n53892), .C(data_tx[2]), .Z(n52582)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;
    defparam n34957_bdd_4_lut_4_lut_else_4_lut.init = 16'h7070;
    FD1P3AX VL53L1X_firm_rdy_i0_i5 (.D(\VL53L1X_data_rx_reg[2] [5]), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(next_VL53L1X_firm_rdy[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_firm_rdy_i0_i5.GSR = "ENABLED";
    FD1P3AX VL53L1X_firm_rdy_i0_i4 (.D(\VL53L1X_data_rx_reg[2] [4]), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(next_VL53L1X_firm_rdy[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_firm_rdy_i0_i4.GSR = "ENABLED";
    FD1P3IX cal_reg_addr_i7 (.D(n47981), .SP(sys_clk_enable_73), .CD(n53891), 
            .CK(sys_clk), .Q(cal_reg_addr[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam cal_reg_addr_i7.GSR = "ENABLED";
    FD1P3AX VL53L1X_firm_rdy_i0_i3 (.D(\VL53L1X_data_rx_reg[2] [3]), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(next_VL53L1X_firm_rdy[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_firm_rdy_i0_i3.GSR = "ENABLED";
    FD1P3AX VL53L1X_firm_rdy_i0_i2 (.D(\VL53L1X_data_rx_reg[2] [2]), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(next_VL53L1X_firm_rdy[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_firm_rdy_i0_i2.GSR = "ENABLED";
    LUT4 i23385_4_lut_4_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n53892), .C(\next_i2c_device_driver_state[2] ), .D(n34032), 
         .Z(n14_adj_5272)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A !(B (C)+!B !(C+!(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam i23385_4_lut_4_lut_4_lut.init = 16'h4340;
    FD1P3AX VL53L1X_firm_rdy_i0_i1 (.D(\VL53L1X_data_rx_reg[2] [1]), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(next_VL53L1X_firm_rdy[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_firm_rdy_i0_i1.GSR = "ENABLED";
    FD1P3IX cal_reg_addr_i6 (.D(n47983), .SP(sys_clk_enable_73), .CD(n53891), 
            .CK(sys_clk), .Q(cal_reg_addr[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam cal_reg_addr_i6.GSR = "ENABLED";
    FD1P3JX cal_reg_addr_i5 (.D(n15_adj_5273), .SP(sys_clk_enable_73), .PD(n53891), 
            .CK(sys_clk), .Q(cal_reg_addr[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam cal_reg_addr_i5.GSR = "ENABLED";
    LUT4 n27327_bdd_4_lut_then_4_lut (.A(\next_i2c_device_driver_state[2] ), 
         .B(n53892), .C(\next_i2c_device_driver_state[0] ), .D(\next_i2c_device_driver_state[3] ), 
         .Z(n52592)) /* synthesis lut_function=(!(A+(B (D)+!B !(C+!(D))))) */ ;
    defparam n27327_bdd_4_lut_then_4_lut.init = 16'h1055;
    LUT4 n27327_bdd_4_lut_else_4_lut (.A(\next_i2c_device_driver_state[2] ), 
         .B(n53892), .C(\next_i2c_device_driver_state[0] ), .D(\next_i2c_device_driver_state[3] ), 
         .Z(n52591)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam n27327_bdd_4_lut_else_4_lut.init = 16'h0040;
    FD1P3AX VL53L1X_range_mm_i0_i15 (.D(n52372), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(next_VL53L1X_range_mm[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_range_mm_i0_i15.GSR = "ENABLED";
    FD1P3AX VL53L1X_range_mm_i0_i14 (.D(n52371), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(next_VL53L1X_range_mm[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_range_mm_i0_i14.GSR = "ENABLED";
    FD1P3AX VL53L1X_range_mm_i0_i13 (.D(n52370), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(next_VL53L1X_range_mm[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_range_mm_i0_i13.GSR = "ENABLED";
    FD1P3AX VL53L1X_data_rdy__i8 (.D(\VL53L1X_data_rx_reg[3] [7]), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(\next_VL53L1X_data_rdy[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_data_rdy__i8.GSR = "ENABLED";
    FD1P3IX cal_reg_addr_i4 (.D(n47982), .SP(sys_clk_enable_73), .CD(n53891), 
            .CK(sys_clk), .Q(cal_reg_addr[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam cal_reg_addr_i4.GSR = "ENABLED";
    FD1P3AX VL53L1X_range_mm_i0_i12 (.D(n52369), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(next_VL53L1X_range_mm[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_range_mm_i0_i12.GSR = "ENABLED";
    FD1P3AX VL53L1X_range_mm_i0_i11 (.D(n52368), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(next_VL53L1X_range_mm[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_range_mm_i0_i11.GSR = "ENABLED";
    FD1P3AX VL53L1X_range_mm_i0_i10 (.D(n52367), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(next_VL53L1X_range_mm[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_range_mm_i0_i10.GSR = "ENABLED";
    FD1P3AX VL53L1X_chip_id_i0_i0 (.D(n52333), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(next_VL53L1X_chip_id[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_chip_id_i0_i0.GSR = "ENABLED";
    FD1P3AX VL53L1X_range_mm_i0_i9 (.D(n52366), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(next_VL53L1X_range_mm[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_range_mm_i0_i9.GSR = "ENABLED";
    FD1P3AX VL53L1X_range_mm_i0_i8 (.D(n52365), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(next_VL53L1X_range_mm[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_range_mm_i0_i8.GSR = "ENABLED";
    FD1P3AX VL53L1X_range_mm_i0_i7 (.D(\VL53L1X_data_rx_reg[7] [7]), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(next_VL53L1X_range_mm[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_range_mm_i0_i7.GSR = "ENABLED";
    LUT4 led_data_out_4__I_0_858_Mux_7_i8_3_lut (.A(cal_reg_addr[7]), .B(data_reg[7]), 
         .C(\next_i2c_device_driver_state[0] ), .Z(n8_adj_5262)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam led_data_out_4__I_0_858_Mux_7_i8_3_lut.init = 16'hcaca;
    FD1P3AX VL53L1X_range_mm_i0_i6 (.D(n52386), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(next_VL53L1X_range_mm[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_range_mm_i0_i6.GSR = "ENABLED";
    FD1P3AX VL53L1X_range_mm_i0_i5 (.D(n52384), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(next_VL53L1X_range_mm[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_range_mm_i0_i5.GSR = "ENABLED";
    FD1P3JX cal_reg_addr_i3 (.D(n15_adj_5274), .SP(sys_clk_enable_73), .PD(n53891), 
            .CK(sys_clk), .Q(cal_reg_addr[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam cal_reg_addr_i3.GSR = "ENABLED";
    FD1P3AX VL53L1X_range_mm_i0_i4 (.D(n52381), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(next_VL53L1X_range_mm[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_range_mm_i0_i4.GSR = "ENABLED";
    FD1P3AX VL53L1X_range_mm_i0_i3 (.D(n52380), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(next_VL53L1X_range_mm[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_range_mm_i0_i3.GSR = "ENABLED";
    FD1P3AX VL53L1X_range_mm_i0_i2 (.D(n52377), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(next_VL53L1X_range_mm[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_range_mm_i0_i2.GSR = "ENABLED";
    FD1P3AX VL53L1X_range_mm_i0_i1 (.D(n52376), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(next_VL53L1X_range_mm[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_range_mm_i0_i1.GSR = "ENABLED";
    FD1P3AX VL53L1X_data_rdy__i7 (.D(\VL53L1X_data_rx_reg[3] [6]), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(\next_VL53L1X_data_rdy[6] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_data_rdy__i7.GSR = "ENABLED";
    FD1P3JX cal_reg_addr_i2 (.D(n15_adj_5275), .SP(sys_clk_enable_73), .PD(n53891), 
            .CK(sys_clk), .Q(cal_reg_addr[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam cal_reg_addr_i2.GSR = "ENABLED";
    FD1P3IX cal_reg_addr_i1 (.D(n47980), .SP(sys_clk_enable_73), .CD(n53891), 
            .CK(sys_clk), .Q(cal_reg_addr[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam cal_reg_addr_i1.GSR = "ENABLED";
    LUT4 i23388_4_lut (.A(n34018), .B(data_reg[1]), .C(\i2c_top_debug[1] ), 
         .D(n27301), .Z(n10_adj_5276)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(53[22:35])
    defparam i23388_4_lut.init = 16'hca0a;
    LUT4 led_data_out_4__I_0_858_Mux_2_i8_3_lut (.A(cal_reg_addr[2]), .B(data_reg[2]), 
         .C(\next_i2c_device_driver_state[0] ), .Z(n8_adj_5263)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam led_data_out_4__I_0_858_Mux_2_i8_3_lut.init = 16'hcaca;
    LUT4 i39950_2_lut_rep_537 (.A(resetn), .B(wd_event_active), .C(n52306), 
         .D(\i2c_top_debug[1] ), .Z(n53891)) /* synthesis lut_function=((B+!(C+(D)))+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(371[14:35])
    defparam i39950_2_lut_rep_537.init = 16'hdddf;
    LUT4 i39765_3_lut_4_lut (.A(n53892), .B(n52246), .C(measurement_period_tx_index[0]), 
         .D(measurement_period_tx_index[1]), .Z(next_measurement_period_tx_index[1])) /* synthesis lut_function=(((C (D)+!C !(D))+!B)+!A) */ ;
    defparam i39765_3_lut_4_lut.init = 16'hf77f;
    FD1P3AX VL53L1X_data_rdy__i6 (.D(\VL53L1X_data_rx_reg[3] [5]), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(\next_VL53L1X_data_rdy[5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_data_rdy__i6.GSR = "ENABLED";
    FD1P3AX VL53L1X_data_rdy__i5 (.D(\VL53L1X_data_rx_reg[3] [4]), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(\next_VL53L1X_data_rdy[4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_data_rdy__i5.GSR = "ENABLED";
    FD1P3AX VL53L1X_data_rdy__i4 (.D(\VL53L1X_data_rx_reg[3] [3]), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(\next_VL53L1X_data_rdy[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_data_rdy__i4.GSR = "ENABLED";
    FD1P3AX VL53L1X_data_rdy__i3 (.D(\VL53L1X_data_rx_reg[3] [2]), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(\next_VL53L1X_data_rdy[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_data_rdy__i3.GSR = "ENABLED";
    FD1S3AY measurement_period_tx_index_i2 (.D(next_measurement_period_tx_index[2]), 
            .CK(sys_clk), .Q(measurement_period_tx_index[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam measurement_period_tx_index_i2.GSR = "ENABLED";
    FD1P3AX VL53L1X_data_rdy__i2 (.D(\VL53L1X_data_rx_reg[3] [1]), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(\next_VL53L1X_data_rdy[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_data_rdy__i2.GSR = "ENABLED";
    PFUMX i38619 (.BLUT(n7_adj_5265), .ALUT(n14_adj_5277), .C0(\next_i2c_device_driver_state[3] ), 
          .Z(n49414));
    LUT4 i66_4_lut (.A(n34018), .B(data_reg[6]), .C(\i2c_top_debug[1] ), 
         .D(n27301), .Z(n24)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(53[22:35])
    defparam i66_4_lut.init = 16'hca0a;
    LUT4 i2_2_lut_rep_504 (.A(n53892), .B(\next_i2c_device_driver_state[0] ), 
         .Z(n52440)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i2_2_lut_rep_504.init = 16'h4444;
    LUT4 i1_3_lut_4_lut (.A(n53892), .B(\next_i2c_device_driver_state[0] ), 
         .C(\next_i2c_device_driver_return_state[0] ), .D(next_i2c_state_4__N_1050[0]), 
         .Z(n37)) /* synthesis lut_function=(!(A+!(B (C+!(D))))) */ ;
    defparam i1_3_lut_4_lut.init = 16'h4044;
    LUT4 n52573_bdd_4_lut (.A(n52573), .B(n52574), .C(\next_i2c_device_driver_state[3] ), 
         .D(\next_i2c_device_driver_state[2] ), .Z(n53879)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n52573_bdd_4_lut.init = 16'h00ca;
    LUT4 i7280_3_lut_rep_291_4_lut (.A(cal_reg_addr[0]), .B(n52403), .C(n27913), 
         .D(cal_reg_addr[7]), .Z(n52227)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (C (D))) */ ;
    defparam i7280_3_lut_rep_291_4_lut.init = 16'hf800;
    LUT4 i27105_4_lut (.A(n21_adj_5269), .B(\next_i2c_device_driver_state[2] ), 
         .C(n28), .D(\next_i2c_device_driver_state[3] ), .Z(n21563)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam i27105_4_lut.init = 16'hc088;
    LUT4 mux_3485_i3_4_lut (.A(n53), .B(\next_i2c_device_driver_state[3] ), 
         .C(n6972), .D(VL53L1X_data_rx_reg_index[2]), .Z(n6915[2])) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(395[14] 871[12])
    defparam mux_3485_i3_4_lut.init = 16'h3530;
    LUT4 i39569_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52336), 
         .Z(VL53L1X_data_rx_reg_1__3__N_708)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39569_3_lut.init = 16'h5757;
    LUT4 i39458_2_lut_3_lut_4_lut (.A(n6974), .B(n52448), .C(n6915[0]), 
         .D(n48780), .Z(VL53L1X_data_rx_reg_index_5__N_463)) /* synthesis lut_function=(A (B+!(D))+!A (B+!(C+(D)))) */ ;
    defparam i39458_2_lut_3_lut_4_lut.init = 16'hccef;
    LUT4 i4_4_lut_adj_317 (.A(n6), .B(n52296), .C(n7250), .D(n49365), 
         .Z(n48780)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;
    defparam i4_4_lut_adj_317.init = 16'hfeff;
    LUT4 i39812_2_lut (.A(\next_i2c_device_driver_state[3] ), .B(\next_i2c_device_driver_state[2] ), 
         .Z(n49547)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i39812_2_lut.init = 16'hdddd;
    CCU2D add_3739_11 (.A0(count_sys_clk_for_ms[9]), .B0(n14126), .C0(GND_net), 
          .D0(GND_net), .A1(count_sys_clk_for_ms[10]), .B1(n14126), .C1(GND_net), 
          .D1(GND_net), .CIN(n43791), .COUT(n43792), .S0(count_sys_clk_for_ms_16__N_874[9]), 
          .S1(count_sys_clk_for_ms_16__N_874[10]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(211[14] 219[12])
    defparam add_3739_11.INIT0 = 16'h7777;
    defparam add_3739_11.INIT1 = 16'h4444;
    defparam add_3739_11.INJECT1_0 = "NO";
    defparam add_3739_11.INJECT1_1 = "NO";
    LUT4 i1_4_lut_4_lut_then_4_lut (.A(\next_i2c_device_driver_state[4] ), 
         .B(\next_i2c_device_driver_state[3] ), .C(\next_i2c_device_driver_state[2] ), 
         .D(n53892), .Z(n52487)) /* synthesis lut_function=(!(A+!(B (D)+!B (C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam i1_4_lut_4_lut_then_4_lut.init = 16'h5410;
    LUT4 n51720_bdd_3_lut (.A(n51720), .B(n46979), .C(\next_i2c_device_driver_state[3] ), 
         .Z(n51721)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n51720_bdd_3_lut.init = 16'hcaca;
    LUT4 i39706_2_lut (.A(\next_i2c_device_driver_state[4] ), .B(\next_i2c_device_driver_state[3] ), 
         .Z(n49665)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i39706_2_lut.init = 16'hbbbb;
    LUT4 n33840_bdd_3_lut_40798 (.A(n33840), .B(n46603), .C(\next_i2c_device_driver_state[3] ), 
         .Z(n51722)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n33840_bdd_3_lut_40798.init = 16'hcaca;
    LUT4 n6_bdd_4_lut (.A(n6), .B(n7246), .C(n52296), .D(\next_i2c_device_driver_state[2] ), 
         .Z(n51725)) /* synthesis lut_function=(A (B (C (D)))+!A (B ((D)+!C))) */ ;
    defparam n6_bdd_4_lut.init = 16'hc404;
    LUT4 i4_4_lut_adj_318 (.A(n7_adj_5278), .B(next_addr_7__N_1168), .C(n53892), 
         .D(n52314), .Z(count_ms_15__N_910[4])) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;
    defparam i4_4_lut_adj_318.init = 16'hfffb;
    LUT4 VL53L1X_data_rx_reg_index_5__N_427_I_0_750_2_lut_3_lut_4_lut (.A(n6974), 
         .B(n52448), .C(n6915[0]), .D(n48780), .Z(VL53L1X_data_rx_reg_index_5__N_445)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam VL53L1X_data_rx_reg_index_5__N_427_I_0_750_2_lut_3_lut_4_lut.init = 16'h0010;
    LUT4 i26061_4_lut (.A(n52137), .B(\next_i2c_device_driver_state[2] ), 
         .C(n28_adj_5279), .D(\next_i2c_device_driver_state[3] ), .Z(n22284)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam i26061_4_lut.init = 16'hc088;
    LUT4 led_data_out_4__I_0_860_Mux_2_i15_4_lut (.A(n7_adj_5267), .B(n53892), 
         .C(\next_i2c_device_driver_state[4] ), .D(n52509), .Z(n15_adj_5280)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam led_data_out_4__I_0_860_Mux_2_i15_4_lut.init = 16'hfaca;
    LUT4 i1_3_lut_4_lut_adj_319 (.A(n52248), .B(next_addr_7__N_1168), .C(n48104), 
         .D(n52420), .Z(n29262)) /* synthesis lut_function=(A (B (C (D))+!B (D))+!A (D)) */ ;
    defparam i1_3_lut_4_lut_adj_319.init = 16'hf700;
    LUT4 i1_4_lut_4_lut_else_4_lut (.A(\next_i2c_device_driver_state[4] ), 
         .B(\next_i2c_device_driver_state[3] ), .C(\next_i2c_device_driver_state[2] ), 
         .D(n53892), .Z(n52486)) /* synthesis lut_function=(!(A+!(B (C+(D))+!B (C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam i1_4_lut_4_lut_else_4_lut.init = 16'h5450;
    LUT4 n47394_bdd_3_lut_40735 (.A(n47394), .B(cal_reg_addr[0]), .C(cal_reg_addr[3]), 
         .Z(n50952)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam n47394_bdd_3_lut_40735.init = 16'h2020;
    LUT4 i19683_3_lut_rep_441 (.A(n30354), .B(n30353), .C(n30352), .Z(n52377)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19683_3_lut_rep_441.init = 16'hcaca;
    LUT4 i39950_2_lut_rep_276_3_lut_4_lut (.A(resetn), .B(wd_event_active), 
         .C(n52306), .D(\i2c_top_debug[1] ), .Z(n52212)) /* synthesis lut_function=((B+!(C+(D)))+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(371[14:35])
    defparam i39950_2_lut_rep_276_3_lut_4_lut.init = 16'hdddf;
    LUT4 i1_3_lut_4_lut_adj_320 (.A(n52248), .B(next_addr_7__N_1168), .C(n48104), 
         .D(n52420), .Z(sys_clk_enable_242)) /* synthesis lut_function=(((C (D))+!B)+!A) */ ;
    defparam i1_3_lut_4_lut_adj_320.init = 16'hf777;
    LUT4 n52582_bdd_4_lut (.A(n52582), .B(n52583), .C(\next_i2c_device_driver_state[3] ), 
         .D(\next_i2c_device_driver_state[2] ), .Z(n53876)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n52582_bdd_4_lut.init = 16'h00ca;
    LUT4 i1_3_lut_4_lut_adj_321 (.A(n52248), .B(next_addr_7__N_1168), .C(n48104), 
         .D(n52449), .Z(sys_clk_enable_255)) /* synthesis lut_function=(((C (D))+!B)+!A) */ ;
    defparam i1_3_lut_4_lut_adj_321.init = 16'hf777;
    LUT4 gnd_bdd_2_lut_40141 (.A(n50950), .B(cal_reg_addr[4]), .Z(n50951)) /* synthesis lut_function=(A (B)) */ ;
    defparam gnd_bdd_2_lut_40141.init = 16'h8888;
    LUT4 i39245_3_lut (.A(n52503), .B(n52506), .C(cal_reg_addr[5]), .Z(n126)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam i39245_3_lut.init = 16'hcaca;
    LUT4 i38934_4_lut_4_lut_4_lut_4_lut (.A(n53892), .B(\next_i2c_device_driver_state[0] ), 
         .C(\next_i2c_device_driver_state[2] ), .D(data_reg[2]), .Z(n49729)) /* synthesis lut_function=(A (C)+!A (((D)+!C)+!B)) */ ;
    defparam i38934_4_lut_4_lut_4_lut_4_lut.init = 16'hf5b5;
    LUT4 cal_reg_addr_1__bdd_4_lut (.A(cal_reg_addr[1]), .B(cal_reg_addr[0]), 
         .C(cal_reg_addr[2]), .D(cal_reg_addr[3]), .Z(n50950)) /* synthesis lut_function=(A (B (C (D)))+!A !(B+(C (D)+!C !(D)))) */ ;
    defparam cal_reg_addr_1__bdd_4_lut.init = 16'h8110;
    LUT4 i1_4_lut (.A(\next_i2c_device_driver_state[2] ), .B(n52154), .C(n19_adj_5281), 
         .D(\next_i2c_device_driver_state[3] ), .Z(n28_adj_5282)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i1_4_lut.init = 16'ha088;
    LUT4 i33210_2_lut (.A(VL53L1X_osc_cal_val[0]), .B(VL53L1X_osc_cal_val[6]), 
         .Z(n2[6])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i33210_2_lut.init = 16'h6666;
    LUT4 i19944_3_lut (.A(n30615), .B(n30614), .C(n30613), .Z(VL53L1X_data_rx_reg_index[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(229[14] 230[75])
    defparam i19944_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_322 (.A(\next_i2c_device_driver_state[2] ), .B(n24_adj_5283), 
         .C(n19_adj_5284), .D(\next_i2c_device_driver_state[3] ), .Z(n28_adj_5285)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i1_4_lut_adj_322.init = 16'ha088;
    FD1S3IX count_sys_clk_for_ms_i16 (.D(count_sys_clk_for_ms_16__N_874[16]), 
            .CK(sys_clk_N_413), .CD(n52172), .Q(count_sys_clk_for_ms[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam count_sys_clk_for_ms_i16.GSR = "ENABLED";
    FD1S3JX count_sys_clk_for_ms_i15 (.D(count_sys_clk_for_ms_16__N_874[15]), 
            .CK(sys_clk_N_413), .PD(n52172), .Q(count_sys_clk_for_ms[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam count_sys_clk_for_ms_i15.GSR = "ENABLED";
    FD1S3IX count_sys_clk_for_ms_i14 (.D(count_sys_clk_for_ms_16__N_874[14]), 
            .CK(sys_clk_N_413), .CD(n52172), .Q(count_sys_clk_for_ms[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam count_sys_clk_for_ms_i14.GSR = "ENABLED";
    FD1S3IX count_sys_clk_for_ms_i13 (.D(count_sys_clk_for_ms_16__N_874[13]), 
            .CK(sys_clk_N_413), .CD(n52172), .Q(count_sys_clk_for_ms[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam count_sys_clk_for_ms_i13.GSR = "ENABLED";
    FD1S3JX count_sys_clk_for_ms_i12 (.D(count_sys_clk_for_ms_16__N_874[12]), 
            .CK(sys_clk_N_413), .PD(n52172), .Q(count_sys_clk_for_ms[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam count_sys_clk_for_ms_i12.GSR = "ENABLED";
    FD1S3IX count_sys_clk_for_ms_i11 (.D(count_sys_clk_for_ms_16__N_874[11]), 
            .CK(sys_clk_N_413), .CD(n52172), .Q(count_sys_clk_for_ms[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam count_sys_clk_for_ms_i11.GSR = "ENABLED";
    FD1S3JX count_sys_clk_for_ms_i10 (.D(count_sys_clk_for_ms_16__N_874[10]), 
            .CK(sys_clk_N_413), .PD(n52172), .Q(count_sys_clk_for_ms[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam count_sys_clk_for_ms_i10.GSR = "ENABLED";
    FD1S3IX count_sys_clk_for_ms_i9 (.D(count_sys_clk_for_ms_16__N_874[9]), 
            .CK(sys_clk_N_413), .CD(n52172), .Q(count_sys_clk_for_ms[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam count_sys_clk_for_ms_i9.GSR = "ENABLED";
    FD1S3IX count_sys_clk_for_ms_i8 (.D(count_sys_clk_for_ms_16__N_874[8]), 
            .CK(sys_clk_N_413), .CD(n52172), .Q(count_sys_clk_for_ms[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam count_sys_clk_for_ms_i8.GSR = "ENABLED";
    FD1S3IX count_sys_clk_for_ms_i7 (.D(count_sys_clk_for_ms_16__N_874[7]), 
            .CK(sys_clk_N_413), .CD(n52172), .Q(count_sys_clk_for_ms[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam count_sys_clk_for_ms_i7.GSR = "ENABLED";
    FD1S3JX count_sys_clk_for_ms_i6 (.D(count_sys_clk_for_ms_16__N_874[6]), 
            .CK(sys_clk_N_413), .PD(n52172), .Q(count_sys_clk_for_ms[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam count_sys_clk_for_ms_i6.GSR = "ENABLED";
    FD1S3JX count_sys_clk_for_ms_i5 (.D(count_sys_clk_for_ms_16__N_874[5]), 
            .CK(sys_clk_N_413), .PD(n52172), .Q(count_sys_clk_for_ms[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam count_sys_clk_for_ms_i5.GSR = "ENABLED";
    FD1S3IX count_sys_clk_for_ms_i4 (.D(count_sys_clk_for_ms_16__N_874[4]), 
            .CK(sys_clk_N_413), .CD(n52172), .Q(count_sys_clk_for_ms[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam count_sys_clk_for_ms_i4.GSR = "ENABLED";
    FD1S3JX count_sys_clk_for_ms_i3 (.D(count_sys_clk_for_ms_16__N_874[3]), 
            .CK(sys_clk_N_413), .PD(n52172), .Q(count_sys_clk_for_ms[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam count_sys_clk_for_ms_i3.GSR = "ENABLED";
    FD1S3JX count_sys_clk_for_ms_i2 (.D(count_sys_clk_for_ms_16__N_874[2]), 
            .CK(sys_clk_N_413), .PD(n52172), .Q(count_sys_clk_for_ms[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam count_sys_clk_for_ms_i2.GSR = "ENABLED";
    LUT4 n6_bdd_2_lut_40691 (.A(n6), .B(n52296), .Z(n51817)) /* synthesis lut_function=((B)+!A) */ ;
    defparam n6_bdd_2_lut_40691.init = 16'hdddd;
    FD1S3JX count_sys_clk_for_ms_i1 (.D(count_sys_clk_for_ms_16__N_874[1]), 
            .CK(sys_clk_N_413), .PD(n52172), .Q(count_sys_clk_for_ms[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam count_sys_clk_for_ms_i1.GSR = "ENABLED";
    FD1S3IX target_read_count_i1 (.D(next_target_read_count_5__N_414[1]), 
            .CK(sys_clk), .CD(n53891), .Q(target_read_count[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam target_read_count_i1.GSR = "ENABLED";
    LUT4 i39221_3_lut_4_lut (.A(cal_reg_addr[3]), .B(n52274), .C(cal_reg_addr[4]), 
         .D(n109), .Z(n125)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;
    defparam i39221_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_5288_i3_4_lut (.A(\next_i2c_device_driver_state[3] ), .B(n52449), 
         .C(n52303), .D(n7244), .Z(n13173[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam mux_5288_i3_4_lut.init = 16'hcacf;
    LUT4 n6_bdd_3_lut_3_lut_4_lut (.A(n53892), .B(\next_i2c_device_driver_state[0] ), 
         .C(\next_i2c_device_driver_return_state[4] ), .D(\next_i2c_device_driver_state[2] ), 
         .Z(n51006)) /* synthesis lut_function=(A+((C+!(D))+!B)) */ ;
    defparam n6_bdd_3_lut_3_lut_4_lut.init = 16'hfbff;
    LUT4 i38716_4_lut_4_lut (.A(n52449), .B(n33834), .C(\next_i2c_device_driver_state[2] ), 
         .D(n37), .Z(n49511)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (B+((D)+!C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i38716_4_lut_4_lut.init = 16'hf5c5;
    LUT4 led_data_out_4__I_0_860_Mux_0_i3_4_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n52270), .C(\next_i2c_device_driver_state[2] ), .D(n69), .Z(n3)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam led_data_out_4__I_0_860_Mux_0_i3_4_lut.init = 16'hcfca;
    LUT4 i17673_2_lut_3_lut (.A(n53892), .B(\next_i2c_device_driver_state[0] ), 
         .C(\next_i2c_device_driver_state[3] ), .Z(n28226)) /* synthesis lut_function=(A (C)+!A (B+(C))) */ ;
    defparam i17673_2_lut_3_lut.init = 16'hf4f4;
    LUT4 i1_2_lut_rep_310_3_lut (.A(resetn), .B(wd_event_active), .C(resetn_imu_N_1182), 
         .Z(n52246)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(371[14:35])
    defparam i1_2_lut_rep_310_3_lut.init = 16'h2020;
    LUT4 i39274_3_lut (.A(n10_adj_5286), .B(n13_adj_5287), .C(\next_i2c_device_driver_state[2] ), 
         .Z(n14_adj_5288)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam i39274_3_lut.init = 16'hcaca;
    CCU2D add_3739_9 (.A0(count_sys_clk_for_ms[7]), .B0(n14126), .C0(GND_net), 
          .D0(GND_net), .A1(count_sys_clk_for_ms[8]), .B1(n14126), .C1(GND_net), 
          .D1(GND_net), .CIN(n43790), .COUT(n43791), .S0(count_sys_clk_for_ms_16__N_874[7]), 
          .S1(count_sys_clk_for_ms_16__N_874[8]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(211[14] 219[12])
    defparam add_3739_9.INIT0 = 16'h7777;
    defparam add_3739_9.INIT1 = 16'h7777;
    defparam add_3739_9.INJECT1_0 = "NO";
    defparam add_3739_9.INJECT1_1 = "NO";
    PFUMX i40932 (.BLUT(n52507), .ALUT(n52508), .C0(\next_i2c_device_driver_state[2] ), 
          .Z(n52509));
    LUT4 i39779_2_lut (.A(n53892), .B(\next_i2c_device_driver_state[3] ), 
         .Z(n30)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i39779_2_lut.init = 16'hbbbb;
    LUT4 i1_2_lut_4_lut (.A(n30354), .B(n30353), .C(n30352), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_7__2__N_504)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut.init = 16'hca00;
    LUT4 mux_3485_i2_4_lut (.A(n53), .B(\next_i2c_device_driver_state[3] ), 
         .C(n6972), .D(n52446), .Z(n6915[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(395[14] 871[12])
    defparam mux_3485_i2_4_lut.init = 16'hcfca;
    LUT4 i1_3_lut_4_lut_adj_323 (.A(n53892), .B(\next_i2c_device_driver_state[0] ), 
         .C(\next_i2c_device_driver_return_state[3] ), .D(next_i2c_state_4__N_1050[0]), 
         .Z(n38)) /* synthesis lut_function=(!(A+!(B (C+!(D))))) */ ;
    defparam i1_3_lut_4_lut_adj_323.init = 16'h4044;
    LUT4 n52579_bdd_4_lut (.A(n52579), .B(n52580), .C(\next_i2c_device_driver_state[3] ), 
         .D(\next_i2c_device_driver_state[2] ), .Z(n53877)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n52579_bdd_4_lut.init = 16'h00ca;
    LUT4 i39858_2_lut_3_lut_4_lut (.A(VL53L1X_data_rx_reg_index[2]), .B(n52444), 
         .C(n52446), .D(n52447), .Z(sys_clk_enable_17)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i39858_2_lut_3_lut_4_lut.init = 16'h0040;
    LUT4 i39896_2_lut_3_lut_4_lut (.A(n52447), .B(n52446), .C(n52444), 
         .D(VL53L1X_data_rx_reg_index[2]), .Z(sys_clk_enable_9)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(229[14] 230[75])
    defparam i39896_2_lut_3_lut_4_lut.init = 16'h0080;
    LUT4 VL53L1X_data_rx_reg_index_i1_i3_3_lut_4_lut (.A(n52447), .B(n52446), 
         .C(one_byte_ready), .D(VL53L1X_data_rx_reg_index[2]), .Z(n23[2])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(229[14] 230[75])
    defparam VL53L1X_data_rx_reg_index_i1_i3_3_lut_4_lut.init = 16'h7f80;
    LUT4 i2_3_lut_4_lut (.A(n52447), .B(n52446), .C(VL53L1X_data_rx_reg_index[2]), 
         .D(n52444), .Z(n28247)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(229[14] 230[75])
    defparam i2_3_lut_4_lut.init = 16'h8000;
    L6MUX21 i38657 (.D0(n49450), .D1(n52136), .SD(\next_i2c_device_driver_state[4] ), 
            .Z(next_data_reg_15__N_362[6]));
    LUT4 mux_5289_i4_4_lut (.A(read_write_in), .B(n52296), .C(n7246), 
         .D(n52203), .Z(n13181[3])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam mux_5289_i4_4_lut.init = 16'hc0ca;
    LUT4 i1_2_lut_3_lut (.A(n53892), .B(\next_i2c_device_driver_state[0] ), 
         .C(\next_i2c_device_driver_return_state[1] ), .Z(n10)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut.init = 16'h4040;
    L6MUX21 i38660 (.D0(n49453), .D1(n49454), .SD(\next_i2c_device_driver_state[4] ), 
            .Z(next_data_reg_15__N_362[3]));
    L6MUX21 i38663 (.D0(n49456), .D1(n49457), .SD(\next_i2c_device_driver_state[4] ), 
            .Z(next_data_reg_15__N_362[1]));
    LUT4 i3_4_lut_rep_360 (.A(n49665), .B(\next_i2c_device_driver_state[0] ), 
         .C(n53892), .D(\next_i2c_device_driver_state[2] ), .Z(n52296)) /* synthesis lut_function=(!(A+(B+!(C (D)+!C !(D))))) */ ;
    defparam i3_4_lut_rep_360.init = 16'h1001;
    LUT4 i27538_2_lut_4_lut (.A(n49665), .B(\next_i2c_device_driver_state[0] ), 
         .C(n53892), .D(\next_i2c_device_driver_state[2] ), .Z(n13144[4])) /* synthesis lut_function=(A+(B+!(C (D)))) */ ;
    defparam i27538_2_lut_4_lut.init = 16'hefff;
    LUT4 i39368_3_lut_4_lut (.A(n52199), .B(\next_i2c_device_driver_state[2] ), 
         .C(\next_i2c_device_driver_state[4] ), .D(n7_adj_5290), .Z(n15_adj_5291)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam i39368_3_lut_4_lut.init = 16'h8f80;
    LUT4 i1_2_lut_rep_333_2_lut_3_lut (.A(n53892), .B(\next_i2c_device_driver_state[0] ), 
         .C(\next_i2c_device_driver_state[2] ), .Z(n52269)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i1_2_lut_rep_333_2_lut_3_lut.init = 16'h0404;
    LUT4 count_ms_15__I_0_875_i9_3_lut (.A(count_ms_15__N_910[4]), .B(count_ms_15__N_894[8]), 
         .C(n7654[7]), .Z(count_ms_15__N_396[8])) /* synthesis lut_function=(A (B (C))+!A (B+!(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(194[14] 219[12])
    defparam count_ms_15__I_0_875_i9_3_lut.init = 16'hc5c5;
    CCU2D add_3739_7 (.A0(count_sys_clk_for_ms[5]), .B0(n14126), .C0(GND_net), 
          .D0(GND_net), .A1(count_sys_clk_for_ms[6]), .B1(n14126), .C1(GND_net), 
          .D1(GND_net), .CIN(n43789), .COUT(n43790), .S0(count_sys_clk_for_ms_16__N_874[5]), 
          .S1(count_sys_clk_for_ms_16__N_874[6]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(211[14] 219[12])
    defparam add_3739_7.INIT0 = 16'h4444;
    defparam add_3739_7.INIT1 = 16'h4444;
    defparam add_3739_7.INJECT1_0 = "NO";
    defparam add_3739_7.INJECT1_1 = "NO";
    LUT4 i39572_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52335), 
         .Z(VL53L1X_data_rx_reg_1__2__N_714)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39572_3_lut.init = 16'h5757;
    LUT4 n51197_bdd_4_lut (.A(n51197), .B(n37158), .C(n51199), .D(n53892), 
         .Z(n52152)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A !((D)+!C)) */ ;
    defparam n51197_bdd_4_lut.init = 16'h88f0;
    LUT4 i11612_3_lut_4_lut (.A(n52292), .B(n52256), .C(data_rx[0]), .D(n52365), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[48])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(252[13:59])
    defparam i11612_3_lut_4_lut.init = 16'hfb40;
    LUT4 i11610_3_lut_4_lut (.A(n52292), .B(n52256), .C(data_rx[1]), .D(n52366), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[49])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(252[13:59])
    defparam i11610_3_lut_4_lut.init = 16'hfb40;
    LUT4 n66_bdd_4_lut_41424 (.A(n66), .B(\next_i2c_device_driver_state[0] ), 
         .C(n52205), .D(next_i2c_state_4__N_1050[0]), .Z(n53051)) /* synthesis lut_function=(A (B+(D))+!A !(B (C)+!B !(D))) */ ;
    defparam n66_bdd_4_lut_41424.init = 16'hbf8c;
    LUT4 i11608_3_lut_4_lut (.A(n52292), .B(n52256), .C(data_rx[2]), .D(n52367), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[50])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(252[13:59])
    defparam i11608_3_lut_4_lut.init = 16'hfb40;
    L6MUX21 i38931 (.D0(n49724), .D1(n49725), .SD(\next_i2c_device_driver_state[4] ), 
            .Z(next_data_reg_15__N_362[7]));
    LUT4 i11606_3_lut_4_lut (.A(n52292), .B(n52256), .C(data_rx[3]), .D(n52368), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[51])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(252[13:59])
    defparam i11606_3_lut_4_lut.init = 16'hfb40;
    L6MUX21 i38938 (.D0(n49731), .D1(n49732), .SD(\next_i2c_device_driver_state[4] ), 
            .Z(next_data_reg_15__N_362[2]));
    LUT4 i11600_3_lut_4_lut (.A(n52292), .B(n52256), .C(data_rx[4]), .D(n52369), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[52])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(252[13:59])
    defparam i11600_3_lut_4_lut.init = 16'hfb40;
    LUT4 n51131_bdd_4_lut (.A(n51131), .B(n37158), .C(n51133), .D(n53892), 
         .Z(n52153)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A !((D)+!C)) */ ;
    defparam n51131_bdd_4_lut.init = 16'h88f0;
    LUT4 n33838_bdd_4_lut_40681 (.A(next_data_tx_7__N_1032[0]), .B(n37517), 
         .C(data_tx[0]), .D(\next_i2c_device_driver_state[0] ), .Z(n51024)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam n33838_bdd_4_lut_40681.init = 16'hc088;
    LUT4 n66_bdd_2_lut_41425 (.A(\next_i2c_state_4__N_1055[1] ), .B(\next_i2c_device_driver_state[0] ), 
         .Z(n53052)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam n66_bdd_2_lut_41425.init = 16'h4444;
    LUT4 i11575_3_lut_4_lut (.A(n52292), .B(n52256), .C(data_rx[5]), .D(n52370), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[53])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(252[13:59])
    defparam i11575_3_lut_4_lut.init = 16'hfb40;
    LUT4 i1_2_lut_4_lut_adj_324 (.A(n30406), .B(n30405), .C(n30404), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_5__5__N_582)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_324.init = 16'hca00;
    LUT4 i11548_3_lut_4_lut (.A(n52292), .B(n52256), .C(data_rx[6]), .D(n52371), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[54])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(252[13:59])
    defparam i11548_3_lut_4_lut.init = 16'hfb40;
    LUT4 i11444_3_lut_4_lut (.A(n52292), .B(n52256), .C(data_rx[7]), .D(n52372), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[55])) /* synthesis lut_function=(A (D)+!A (B (C)+!B (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(252[13:59])
    defparam i11444_3_lut_4_lut.init = 16'hfb40;
    LUT4 n6_bdd_3_lut_3_lut_4_lut_adj_325 (.A(\next_i2c_device_driver_state[2] ), 
         .B(n52460), .C(next_imu_good), .D(n52449), .Z(n51724)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;
    defparam n6_bdd_3_lut_3_lut_4_lut_adj_325.init = 16'hf7ff;
    LUT4 i26993_2_lut_3_lut_4_lut (.A(\next_i2c_device_driver_state[2] ), 
         .B(n52460), .C(read_write_in), .D(sys_clk_enable_108), .Z(n13173[1])) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (C+!(D))) */ ;
    defparam i26993_2_lut_3_lut_4_lut.init = 16'hf0f7;
    LUT4 i10059_3_lut_4_lut (.A(\next_i2c_device_driver_state[2] ), .B(n52460), 
         .C(n53892), .D(n7244), .Z(n20052)) /* synthesis lut_function=(!(A (B (C)+!B (D))+!A (D))) */ ;
    defparam i10059_3_lut_4_lut.init = 16'h087f;
    LUT4 i27029_4_lut (.A(n52153), .B(\next_i2c_device_driver_state[2] ), 
         .C(n28_adj_5292), .D(\next_i2c_device_driver_state[3] ), .Z(n23389)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam i27029_4_lut.init = 16'hc088;
    LUT4 n51101_bdd_4_lut (.A(n51101), .B(n37158), .C(n51103), .D(n53892), 
         .Z(n52154)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A !((D)+!C)) */ ;
    defparam n51101_bdd_4_lut.init = 16'h88f0;
    LUT4 next_i2c_device_driver_state_1__bdd_4_lut_41238 (.A(\next_i2c_device_driver_state[2] ), 
         .B(\next_i2c_state_4__N_1055[1] ), .C(\next_i2c_device_driver_state[0] ), 
         .D(n72), .Z(n53050)) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C+(D)))) */ ;
    defparam next_i2c_device_driver_state_1__bdd_4_lut_41238.init = 16'hff10;
    LUT4 measurement_period_tx_index_0__bdd_3_lut (.A(VL53L1X_measurement_period[0]), 
         .B(measurement_period_tx_index[1]), .C(VL53L1X_measurement_period[16]), 
         .Z(n52077)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam measurement_period_tx_index_0__bdd_3_lut.init = 16'he2e2;
    LUT4 measurement_period_tx_index_0__bdd_2_lut (.A(measurement_period_tx_index[1]), 
         .B(VL53L1X_measurement_period[8]), .Z(n52076)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam measurement_period_tx_index_0__bdd_2_lut.init = 16'h4444;
    LUT4 i25867_2_lut_rep_378 (.A(\next_i2c_device_driver_state[2] ), .B(\next_i2c_device_driver_state[3] ), 
         .Z(n52314)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam i25867_2_lut_rep_378.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_adj_326 (.A(\next_i2c_device_driver_state[2] ), .B(\next_i2c_device_driver_state[3] ), 
         .C(\next_i2c_device_driver_state[4] ), .Z(n49226)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam i1_2_lut_3_lut_adj_326.init = 16'hfefe;
    LUT4 n52087_bdd_3_lut (.A(n52087), .B(n52085), .C(\next_i2c_device_driver_state[4] ), 
         .Z(next_i2c_state_4__N_386[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n52087_bdd_3_lut.init = 16'hcaca;
    LUT4 i39801_2_lut (.A(\next_i2c_device_driver_state[2] ), .B(n53892), 
         .Z(n37517)) /* synthesis lut_function=(!(A+(B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i39801_2_lut.init = 16'h1111;
    LUT4 n6_bdd_4_lut_adj_327 (.A(\next_i2c_device_driver_state[0] ), .B(\next_i2c_device_driver_return_state[4] ), 
         .C(next_i2c_state_4__N_1050[0]), .D(n53892), .Z(n52122)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (D)) */ ;
    defparam n6_bdd_4_lut_adj_327.init = 16'hff80;
    CCU2D add_3739_5 (.A0(count_sys_clk_for_ms[3]), .B0(n14126), .C0(GND_net), 
          .D0(GND_net), .A1(count_sys_clk_for_ms[4]), .B1(n14126), .C1(GND_net), 
          .D1(GND_net), .CIN(n43788), .COUT(n43789), .S0(count_sys_clk_for_ms_16__N_874[3]), 
          .S1(count_sys_clk_for_ms_16__N_874[4]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(211[14] 219[12])
    defparam add_3739_5.INIT0 = 16'h4444;
    defparam add_3739_5.INIT1 = 16'h7777;
    defparam add_3739_5.INJECT1_0 = "NO";
    defparam add_3739_5.INJECT1_1 = "NO";
    PFUMX i38661 (.BLUT(n7_adj_5293), .ALUT(n14_adj_5272), .C0(\next_i2c_device_driver_state[3] ), 
          .Z(n49456));
    PFUMX i38658 (.BLUT(n7_adj_5294), .ALUT(n14_adj_5295), .C0(\next_i2c_device_driver_state[3] ), 
          .Z(n49453));
    PFUMX i38655 (.BLUT(n7_adj_5264), .ALUT(n14_adj_5296), .C0(\next_i2c_device_driver_state[3] ), 
          .Z(n49450));
    LUT4 i2_3_lut (.A(cal_reg_addr[2]), .B(n27913), .C(cal_reg_addr[1]), 
         .Z(n47344)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut.init = 16'hfefe;
    FD1P3IX VL53L1X_measurement_period__i20 (.D(next_VL53L1X_measurement_period_31__N_1103[22]), 
            .SP(sys_clk_enable_108), .CD(n53891), .CK(sys_clk), .Q(VL53L1X_measurement_period[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam VL53L1X_measurement_period__i20.GSR = "ENABLED";
    PFUMX i40930 (.BLUT(n52504), .ALUT(n52505), .C0(cal_reg_addr[0]), 
          .Z(n52506));
    LUT4 i3_4_lut (.A(cal_reg_addr[3]), .B(cal_reg_addr[6]), .C(cal_reg_addr[4]), 
         .D(cal_reg_addr[5]), .Z(n27913)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i3_4_lut.init = 16'hfffe;
    LUT4 n7_bdd_3_lut (.A(n7_adj_5267), .B(n52123), .C(\next_i2c_device_driver_state[3] ), 
         .Z(n52124)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n7_bdd_3_lut.init = 16'hcaca;
    LUT4 i19675_3_lut_rep_445 (.A(n30346), .B(n30345), .C(n30344), .Z(n52381)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19675_3_lut_rep_445.init = 16'hcaca;
    LUT4 n52576_bdd_4_lut (.A(n52576), .B(n52577), .C(\next_i2c_device_driver_state[3] ), 
         .D(\next_i2c_device_driver_state[2] ), .Z(n53878)) /* synthesis lut_function=(!(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B))) */ ;
    defparam n52576_bdd_4_lut.init = 16'h00ca;
    FD1P3IX VL53L1X_measurement_period__i19 (.D(next_VL53L1X_measurement_period_31__N_1103[21]), 
            .SP(sys_clk_enable_108), .CD(n53891), .CK(sys_clk), .Q(VL53L1X_measurement_period[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam VL53L1X_measurement_period__i19.GSR = "ENABLED";
    LUT4 i1_2_lut_4_lut_adj_328 (.A(n30350), .B(n30349), .C(n30348), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_7__3__N_498)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_328.init = 16'hca00;
    FD1P3IX VL53L1X_measurement_period__i18 (.D(next_VL53L1X_measurement_period_31__N_1103[20]), 
            .SP(sys_clk_enable_108), .CD(n53891), .CK(sys_clk), .Q(VL53L1X_measurement_period[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam VL53L1X_measurement_period__i18.GSR = "ENABLED";
    LUT4 i27134_4_lut (.A(VL53L1X_measurement_period[6]), .B(n52445), .C(VL53L1X_measurement_period[14]), 
         .D(measurement_period_tx_index[0]), .Z(next_data_tx_7__N_1024[6])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(721[21] 727[28])
    defparam i27134_4_lut.init = 16'h3022;
    LUT4 i19679_3_lut_rep_444 (.A(n30350), .B(n30349), .C(n30348), .Z(n52380)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19679_3_lut_rep_444.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_329 (.A(n30346), .B(n30345), .C(n30344), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_7__4__N_492)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_329.init = 16'hca00;
    FD1P3IX VL53L1X_measurement_period__i17 (.D(next_VL53L1X_measurement_period_31__N_1103[19]), 
            .SP(sys_clk_enable_108), .CD(n53891), .CK(sys_clk), .Q(VL53L1X_measurement_period[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam VL53L1X_measurement_period__i17.GSR = "ENABLED";
    LUT4 i19755_3_lut (.A(n30426), .B(n30425), .C(n30424), .Z(\VL53L1X_data_rx_reg[5] [0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19755_3_lut.init = 16'hcaca;
    FD1P3IX VL53L1X_measurement_period__i16 (.D(next_VL53L1X_measurement_period_31__N_1103[18]), 
            .SP(sys_clk_enable_108), .CD(n53891), .CK(sys_clk), .Q(VL53L1X_measurement_period[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam VL53L1X_measurement_period__i16.GSR = "ENABLED";
    LUT4 i19671_3_lut_rep_448 (.A(n30342), .B(n30341), .C(n30340), .Z(n52384)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19671_3_lut_rep_448.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_330 (.A(n30342), .B(n30341), .C(n30340), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_7__5__N_486)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_330.init = 16'hca00;
    LUT4 i19667_3_lut_rep_450 (.A(n30338), .B(n30337), .C(n30336), .Z(n52386)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19667_3_lut_rep_450.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_331 (.A(n30338), .B(n30337), .C(n30336), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_7__6__N_480)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_331.init = 16'hca00;
    FD1P3IX VL53L1X_measurement_period__i15 (.D(next_VL53L1X_measurement_period_31__N_1103[17]), 
            .SP(sys_clk_enable_108), .CD(n53891), .CK(sys_clk), .Q(VL53L1X_measurement_period[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam VL53L1X_measurement_period__i15.GSR = "ENABLED";
    PFUMX i51 (.BLUT(n16), .ALUT(n20_adj_5297), .C0(n53892), .Z(n24_adj_5283));
    LUT4 i1_4_lut_4_lut_adj_332 (.A(next_i2c_state_4__N_1050[0]), .B(n52440), 
         .C(n33834), .D(\next_i2c_device_driver_return_state[2] ), .Z(n13_adj_5287)) /* synthesis lut_function=(A (B (C+(D))+!B (C))+!A (B+(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam i1_4_lut_4_lut_adj_332.init = 16'hfcf4;
    FD1P3IX VL53L1X_measurement_period__i14 (.D(next_VL53L1X_measurement_period_31__N_1103[16]), 
            .SP(sys_clk_enable_108), .CD(n53891), .CK(sys_clk), .Q(VL53L1X_measurement_period[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam VL53L1X_measurement_period__i14.GSR = "ENABLED";
    LUT4 i19851_3_lut_rep_384 (.A(n30522), .B(n30521), .C(n30520), .Z(n52320)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19851_3_lut_rep_384.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_333 (.A(n30522), .B(n30521), .C(n30520), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_0__0__N_772)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_333.init = 16'hca00;
    LUT4 i39792_2_lut (.A(\next_i2c_device_driver_state[4] ), .B(\next_i2c_device_driver_state[3] ), 
         .Z(n49571)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam i39792_2_lut.init = 16'heeee;
    LUT4 i39461_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(\VL53L1X_data_rx_reg[7] [7]), 
         .Z(VL53L1X_data_rx_reg_7__7__N_476)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39461_3_lut.init = 16'h5757;
    LUT4 i19847_3_lut_rep_385 (.A(n30518), .B(n30517), .C(n30516), .Z(n52321)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19847_3_lut_rep_385.init = 16'hcaca;
    LUT4 i19663_3_lut (.A(n30334), .B(n30333), .C(n30332), .Z(\VL53L1X_data_rx_reg[7] [7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19663_3_lut.init = 16'hcaca;
    FD1P3IX VL53L1X_measurement_period__i13 (.D(next_VL53L1X_measurement_period_31__N_1103[15]), 
            .SP(sys_clk_enable_108), .CD(n53891), .CK(sys_clk), .Q(VL53L1X_measurement_period[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam VL53L1X_measurement_period__i13.GSR = "ENABLED";
    LUT4 i1_2_lut_4_lut_adj_334 (.A(n30518), .B(n30517), .C(n30516), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_0__1__N_766)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_334.init = 16'hca00;
    LUT4 i19843_3_lut_rep_386 (.A(n30514), .B(n30513), .C(n30512), .Z(n52322)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19843_3_lut_rep_386.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_335 (.A(n30514), .B(n30513), .C(n30512), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_0__2__N_760)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_335.init = 16'hca00;
    FD1P3IX VL53L1X_measurement_period__i12 (.D(next_VL53L1X_measurement_period_31__N_1103[14]), 
            .SP(sys_clk_enable_108), .CD(n53891), .CK(sys_clk), .Q(VL53L1X_measurement_period[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam VL53L1X_measurement_period__i12.GSR = "ENABLED";
    FD1P3IX VL53L1X_measurement_period__i11 (.D(next_VL53L1X_measurement_period_31__N_1103[13]), 
            .SP(sys_clk_enable_108), .CD(n53891), .CK(sys_clk), .Q(VL53L1X_measurement_period[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam VL53L1X_measurement_period__i11.GSR = "ENABLED";
    FD1P3IX VL53L1X_measurement_period__i10 (.D(next_VL53L1X_measurement_period_31__N_1103[12]), 
            .SP(sys_clk_enable_108), .CD(n53891), .CK(sys_clk), .Q(VL53L1X_measurement_period[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam VL53L1X_measurement_period__i10.GSR = "ENABLED";
    PFUMX i38620 (.BLUT(n22), .ALUT(n29_adj_5298), .C0(\next_i2c_device_driver_state[3] ), 
          .Z(n49415));
    LUT4 VL53L1X_measurement_period_3__bdd_2_lut_40403 (.A(VL53L1X_measurement_period[11]), 
         .B(measurement_period_tx_index[1]), .Z(n51099)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam VL53L1X_measurement_period_3__bdd_2_lut_40403.init = 16'h2222;
    FD1P3IX VL53L1X_measurement_period__i9 (.D(next_VL53L1X_measurement_period_31__N_1103[11]), 
            .SP(sys_clk_enable_108), .CD(n53891), .CK(sys_clk), .Q(VL53L1X_measurement_period[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam VL53L1X_measurement_period__i9.GSR = "ENABLED";
    FD1P3IX VL53L1X_measurement_period__i8 (.D(next_VL53L1X_measurement_period_31__N_1103[10]), 
            .SP(sys_clk_enable_108), .CD(n53891), .CK(sys_clk), .Q(VL53L1X_measurement_period[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam VL53L1X_measurement_period__i8.GSR = "ENABLED";
    LUT4 VL53L1X_measurement_period_3__bdd_3_lut_40404 (.A(VL53L1X_measurement_period[3]), 
         .B(measurement_period_tx_index[1]), .C(VL53L1X_measurement_period[19]), 
         .Z(n51100)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam VL53L1X_measurement_period_3__bdd_3_lut_40404.init = 16'he2e2;
    FD1P3IX VL53L1X_measurement_period__i7 (.D(next_VL53L1X_measurement_period_31__N_1103[9]), 
            .SP(sys_clk_enable_108), .CD(n53891), .CK(sys_clk), .Q(VL53L1X_measurement_period[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam VL53L1X_measurement_period__i7.GSR = "ENABLED";
    CCU2D add_3739_3 (.A0(count_sys_clk_for_ms[1]), .B0(n14126), .C0(GND_net), 
          .D0(GND_net), .A1(count_sys_clk_for_ms[2]), .B1(n14126), .C1(GND_net), 
          .D1(GND_net), .CIN(n43787), .COUT(n43788), .S0(count_sys_clk_for_ms_16__N_874[1]), 
          .S1(count_sys_clk_for_ms_16__N_874[2]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(211[14] 219[12])
    defparam add_3739_3.INIT0 = 16'h4444;
    defparam add_3739_3.INIT1 = 16'h4444;
    defparam add_3739_3.INJECT1_0 = "NO";
    defparam add_3739_3.INJECT1_1 = "NO";
    LUT4 i19839_3_lut_rep_388 (.A(n30510), .B(n30509), .C(n30508), .Z(n52324)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19839_3_lut_rep_388.init = 16'hcaca;
    FD1P3IX VL53L1X_measurement_period__i6 (.D(next_VL53L1X_measurement_period_31__N_1103[8]), 
            .SP(sys_clk_enable_108), .CD(n53891), .CK(sys_clk), .Q(VL53L1X_measurement_period[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam VL53L1X_measurement_period__i6.GSR = "ENABLED";
    FD1P3IX VL53L1X_measurement_period__i5 (.D(next_VL53L1X_measurement_period_31__N_1103[7]), 
            .SP(sys_clk_enable_108), .CD(n53891), .CK(sys_clk), .Q(VL53L1X_measurement_period[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam VL53L1X_measurement_period__i5.GSR = "ENABLED";
    FD1S3IX master_trigger_count_ms_i20 (.D(master_trigger_count_ms_20__N_997[20]), 
            .CK(sys_clk), .CD(n52182), .Q(master_trigger_count_ms[20])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(268[14] 281[12])
    defparam master_trigger_count_ms_i20.GSR = "ENABLED";
    PFUMX i40928 (.BLUT(n52501), .ALUT(n52502), .C0(cal_reg_addr[2]), 
          .Z(n52503));
    CCU2D add_3739_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count_sys_clk_for_ms[16]), .B1(n14054), .C1(count_ms[15]), 
          .D1(count_sys_clk_for_ms[0]), .COUT(n43787), .S1(count_sys_clk_for_ms_16__N_874[0]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(211[14] 219[12])
    defparam add_3739_1.INIT0 = 16'h0000;
    defparam add_3739_1.INIT1 = 16'h55a9;
    defparam add_3739_1.INJECT1_0 = "NO";
    defparam add_3739_1.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_336 (.A(\next_i2c_device_driver_state[0] ), .B(n52318), 
         .C(resetn_imu_N_1182), .D(n66), .Z(n72)) /* synthesis lut_function=(A+!(B+!(C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam i1_4_lut_adj_336.init = 16'hbaaa;
    FD1P3IX master_trigger_count_ms_i18 (.D(n611[18]), .SP(sys_clk_enable_224), 
            .CD(n52182), .CK(sys_clk), .Q(master_trigger_count_ms[18])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(268[14] 281[12])
    defparam master_trigger_count_ms_i18.GSR = "ENABLED";
    LUT4 n37158_bdd_2_lut_40249 (.A(data_tx[3]), .B(\next_i2c_device_driver_state[0] ), 
         .Z(n51103)) /* synthesis lut_function=(A (B)) */ ;
    defparam n37158_bdd_2_lut_40249.init = 16'h8888;
    LUT4 i2_3_lut_4_lut_adj_337 (.A(\i2c_top_debug[1] ), .B(\i2c_top_debug[3] ), 
         .C(\i2c_top_debug[4] ), .D(n53886), .Z(n47760)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(53[22:35])
    defparam i2_3_lut_4_lut_adj_337.init = 16'h8000;
    FD1P3IX master_trigger_count_ms_i14 (.D(n611[14]), .SP(sys_clk_enable_224), 
            .CD(n52182), .CK(sys_clk), .Q(master_trigger_count_ms[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(268[14] 281[12])
    defparam master_trigger_count_ms_i14.GSR = "ENABLED";
    LUT4 i1_2_lut_4_lut_adj_338 (.A(n30510), .B(n30509), .C(n30508), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_0__3__N_754)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_338.init = 16'hca00;
    LUT4 i1_2_lut_3_lut_4_lut (.A(\i2c_top_debug[1] ), .B(\i2c_top_debug[3] ), 
         .C(n52425), .D(n51003), .Z(n48098)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(53[22:35])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0800;
    FD1P3IX master_trigger_count_ms_i13 (.D(n611[13]), .SP(sys_clk_enable_224), 
            .CD(n52182), .CK(sys_clk), .Q(master_trigger_count_ms[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(268[14] 281[12])
    defparam master_trigger_count_ms_i13.GSR = "ENABLED";
    FD1P3IX VL53L1X_measurement_period__i4 (.D(next_VL53L1X_measurement_period_31__N_1103[6]), 
            .SP(sys_clk_enable_108), .CD(n53891), .CK(sys_clk), .Q(VL53L1X_measurement_period[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam VL53L1X_measurement_period__i4.GSR = "ENABLED";
    FD1S3IX data_tx__i0 (.D(next_data_tx_7__N_378[0]), .CK(sys_clk), .CD(n53891), 
            .Q(data_tx[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam data_tx__i0.GSR = "ENABLED";
    PFUMX i41220 (.BLUT(n53055), .ALUT(n53054), .C0(\next_i2c_device_driver_state[3] ), 
          .Z(n53056));
    LUT4 i26502_4_lut (.A(measurement_period_tx_index[2]), .B(n52246), .C(n21_adj_5299), 
         .D(n29262), .Z(next_measurement_period_tx_index[2])) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(395[14] 871[12])
    defparam i26502_4_lut.init = 16'hc088;
    LUT4 i11631_2_lut_rep_467 (.A(cal_reg_addr[1]), .B(cal_reg_addr[2]), 
         .Z(n52403)) /* synthesis lut_function=(A (B)) */ ;
    defparam i11631_2_lut_rep_467.init = 16'h8888;
    LUT4 i26022_2_lut_rep_338_3_lut (.A(cal_reg_addr[1]), .B(cal_reg_addr[2]), 
         .C(cal_reg_addr[0]), .Z(n52274)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i26022_2_lut_rep_338_3_lut.init = 16'h8080;
    LUT4 i2_3_lut_4_lut_adj_339 (.A(cal_reg_addr[1]), .B(cal_reg_addr[2]), 
         .C(cal_reg_addr[5]), .D(cal_reg_addr[4]), .Z(n47394)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2_3_lut_4_lut_adj_339.init = 16'h8000;
    LUT4 i26884_4_lut (.A(measurement_period_tx_index[2]), .B(n53892), .C(measurement_period_tx_index[1]), 
         .D(measurement_period_tx_index[0]), .Z(n21_adj_5299)) /* synthesis lut_function=(A (B (C+(D)))+!A !((C+(D))+!B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam i26884_4_lut.init = 16'h8884;
    FD1P3IX VL53L1X_measurement_period__i3 (.D(next_VL53L1X_measurement_period_31__N_1103[5]), 
            .SP(sys_clk_enable_108), .CD(n53891), .CK(sys_clk), .Q(VL53L1X_measurement_period[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam VL53L1X_measurement_period__i3.GSR = "ENABLED";
    FD1P3IX master_trigger_count_ms_i10 (.D(n611[10]), .SP(sys_clk_enable_224), 
            .CD(n52182), .CK(sys_clk), .Q(master_trigger_count_ms[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(268[14] 281[12])
    defparam master_trigger_count_ms_i10.GSR = "ENABLED";
    FD1P3IX VL53L1X_measurement_period__i2 (.D(next_VL53L1X_measurement_period_31__N_1103[4]), 
            .SP(sys_clk_enable_108), .CD(n53891), .CK(sys_clk), .Q(VL53L1X_measurement_period[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam VL53L1X_measurement_period__i2.GSR = "ENABLED";
    FD1P3IX master_trigger_count_ms_i9 (.D(n611[9]), .SP(sys_clk_enable_224), 
            .CD(n52182), .CK(sys_clk), .Q(master_trigger_count_ms[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(268[14] 281[12])
    defparam master_trigger_count_ms_i9.GSR = "ENABLED";
    LUT4 mux_3602_i3_4_lut (.A(n51819), .B(is_2_byte_reg), .C(n7250), 
         .D(n52231), .Z(n2485[2])) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam mux_3602_i3_4_lut.init = 16'hfaca;
    FD1P3IX VL53L1X_measurement_period__i1 (.D(next_VL53L1X_measurement_period_31__N_1103[3]), 
            .SP(sys_clk_enable_108), .CD(n53891), .CK(sys_clk), .Q(VL53L1X_measurement_period[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam VL53L1X_measurement_period__i1.GSR = "ENABLED";
    CCU2D add_409_3 (.A0(cal_reg_addr[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cal_reg_addr[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43783), .COUT(n43784), .S0(next_cal_reg_addr_7__N_1124[1]), 
          .S1(next_cal_reg_addr_7__N_1124[2]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(602[42:66])
    defparam add_409_3.INIT0 = 16'h5aaa;
    defparam add_409_3.INIT1 = 16'h5aaa;
    defparam add_409_3.INJECT1_0 = "NO";
    defparam add_409_3.INJECT1_1 = "NO";
    LUT4 i39920_4_lut (.A(n52271), .B(\next_i2c_device_driver_state[4] ), 
         .C(\next_i2c_device_driver_state[3] ), .D(n52269), .Z(sys_clk_enable_73)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+!((D)+!C)))) */ ;
    defparam i39920_4_lut.init = 16'h3101;
    LUT4 i38842_2_lut (.A(cal_reg_addr[7]), .B(cal_reg_addr[6]), .Z(n49637)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i38842_2_lut.init = 16'h4444;
    FD1S3IX return_state__i5 (.D(next_return_state_4__N_391[4]), .CK(sys_clk), 
            .CD(n53891), .Q(\next_i2c_device_driver_return_state[4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam return_state__i5.GSR = "ENABLED";
    LUT4 led_data_out_4__I_0_860_Mux_1_i29_4_lut_4_lut (.A(\next_i2c_device_driver_state[3] ), 
         .B(\next_i2c_state_4__N_1055[1] ), .C(n52233), .D(n52440), .Z(n29_adj_5300)) /* synthesis lut_function=(A (B (D))+!A !(C)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam led_data_out_4__I_0_860_Mux_1_i29_4_lut_4_lut.init = 16'h8d05;
    LUT4 i12262_3_lut_4_lut (.A(n52447), .B(n52218), .C(data_rx[0]), .D(\VL53L1X_data_rx_reg[5] [0]), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[40])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(252[13:59])
    defparam i12262_3_lut_4_lut.init = 16'hfd20;
    FD1P3IX master_trigger_count_ms_i8 (.D(n611[8]), .SP(sys_clk_enable_224), 
            .CD(n52182), .CK(sys_clk), .Q(master_trigger_count_ms[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(268[14] 281[12])
    defparam master_trigger_count_ms_i8.GSR = "ENABLED";
    LUT4 led_data_out_4__I_0_868_Mux_0_i15_4_lut (.A(n52271), .B(next_cal_reg_addr_7__N_1124[0]), 
         .C(\next_i2c_device_driver_state[3] ), .D(n52269), .Z(n15)) /* synthesis lut_function=(A (B (C (D)))+!A (B ((D)+!C)+!B !(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam led_data_out_4__I_0_868_Mux_0_i15_4_lut.init = 16'hc505;
    LUT4 i12220_3_lut_4_lut (.A(n52447), .B(n52218), .C(data_rx[1]), .D(n52352), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[41])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(252[13:59])
    defparam i12220_3_lut_4_lut.init = 16'hfd20;
    FD1S3IX return_state__i4 (.D(next_return_state_4__N_391[3]), .CK(sys_clk), 
            .CD(n53891), .Q(\next_i2c_device_driver_return_state[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam return_state__i4.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_340 (.A(\next_i2c_device_driver_state[2] ), .B(n52409), 
         .C(n53892), .D(\next_i2c_device_driver_state[3] ), .Z(n7244)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(B (C (D))))) */ ;
    defparam i1_4_lut_adj_340.init = 16'h4080;
    PFUMX i40926 (.BLUT(n52498), .ALUT(n52499), .C0(\next_i2c_device_driver_state[0] ), 
          .Z(n6));
    FD1S3IX return_state__i3 (.D(next_return_state_4__N_391[2]), .CK(sys_clk), 
            .CD(n53891), .Q(\next_i2c_device_driver_return_state[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam return_state__i3.GSR = "ENABLED";
    FD1S3IX return_state__i2 (.D(next_return_state_4__N_391[1]), .CK(sys_clk), 
            .CD(n53891), .Q(\next_i2c_device_driver_return_state[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam return_state__i2.GSR = "ENABLED";
    LUT4 i3_4_lut_adj_341 (.A(n7_adj_5301), .B(\next_i2c_device_driver_state[3] ), 
         .C(\next_i2c_device_driver_state[0] ), .D(\next_i2c_device_driver_state[4] ), 
         .Z(n7234)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i3_4_lut_adj_341.init = 16'h0020;
    LUT4 i12187_3_lut_4_lut (.A(n52447), .B(n52218), .C(data_rx[2]), .D(n52354), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[42])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(252[13:59])
    defparam i12187_3_lut_4_lut.init = 16'hfd20;
    LUT4 VL53L1X_measurement_period_4__bdd_3_lut_40323 (.A(VL53L1X_measurement_period[4]), 
         .B(measurement_period_tx_index[1]), .C(VL53L1X_measurement_period[20]), 
         .Z(n51130)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam VL53L1X_measurement_period_4__bdd_3_lut_40323.init = 16'he2e2;
    LUT4 i39735_2_lut (.A(\next_i2c_device_driver_state[3] ), .B(\next_i2c_device_driver_state[2] ), 
         .Z(n49625)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i39735_2_lut.init = 16'h7777;
    LUT4 i11636_3_lut_4_lut (.A(n52447), .B(n52218), .C(data_rx[3]), .D(n52357), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[43])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(252[13:59])
    defparam i11636_3_lut_4_lut.init = 16'hfd20;
    LUT4 i11620_3_lut_4_lut (.A(n52447), .B(n52218), .C(data_rx[4]), .D(n52358), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[44])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(252[13:59])
    defparam i11620_3_lut_4_lut.init = 16'hfd20;
    LUT4 i39793_2_lut (.A(\next_i2c_device_driver_state[2] ), .B(n53892), 
         .Z(n49569)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i39793_2_lut.init = 16'heeee;
    LUT4 i11618_3_lut_4_lut (.A(n52447), .B(n52218), .C(data_rx[5]), .D(n52360), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[45])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(252[13:59])
    defparam i11618_3_lut_4_lut.init = 16'hfd20;
    FD1S3IX i2c_state__i5 (.D(next_i2c_state_4__N_386[4]), .CK(sys_clk), 
            .CD(n53891), .Q(\next_i2c_device_driver_state[4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam i2c_state__i5.GSR = "ENABLED";
    LUT4 i1_4_lut_4_lut_else_3_lut_adj_342 (.A(\next_i2c_device_driver_state[3] ), 
         .B(\next_i2c_device_driver_state[0] ), .C(\next_i2c_state_4__N_1055[1] ), 
         .Z(n52507)) /* synthesis lut_function=(!(A ((C)+!B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i1_4_lut_4_lut_else_3_lut_adj_342.init = 16'h5d5d;
    LUT4 i11616_3_lut_4_lut (.A(n52447), .B(n52218), .C(data_rx[6]), .D(n52363), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[46])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(252[13:59])
    defparam i11616_3_lut_4_lut.init = 16'hfd20;
    PFUMX i41218 (.BLUT(n53052), .ALUT(n53051), .C0(\next_i2c_device_driver_state[2] ), 
          .Z(n53053));
    LUT4 i6225_2_lut (.A(count_ms[15]), .B(count_sys_clk_for_ms[16]), .Z(n14126)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(211[14] 219[12])
    defparam i6225_2_lut.init = 16'hbbbb;
    LUT4 i1_2_lut_rep_473 (.A(\next_i2c_device_driver_state[0] ), .B(\next_i2c_device_driver_state[4] ), 
         .Z(n52409)) /* synthesis lut_function=(A (B)) */ ;
    defparam i1_2_lut_rep_473.init = 16'h8888;
    LUT4 VL53L1X_measurement_period_4__bdd_2_lut_40322 (.A(VL53L1X_measurement_period[12]), 
         .B(measurement_period_tx_index[1]), .Z(n51129)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam VL53L1X_measurement_period_4__bdd_2_lut_40322.init = 16'h2222;
    LUT4 i38896_2_lut_rep_474 (.A(\next_i2c_device_driver_state[3] ), .B(\next_i2c_device_driver_state[2] ), 
         .Z(n52410)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i38896_2_lut_rep_474.init = 16'h4444;
    LUT4 i39205_3_lut_4_lut (.A(\next_i2c_device_driver_state[3] ), .B(\next_i2c_device_driver_state[2] ), 
         .C(n52485), .D(n21_adj_5302), .Z(n49478)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;
    defparam i39205_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i1_2_lut_3_lut_adj_343 (.A(\next_i2c_device_driver_state[3] ), .B(\next_i2c_device_driver_state[2] ), 
         .C(\next_i2c_device_driver_state[4] ), .Z(n48104)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;
    defparam i1_2_lut_3_lut_adj_343.init = 16'h4040;
    LUT4 i22_4_lut_4_lut_4_lut_4_lut (.A(\next_i2c_device_driver_state[3] ), 
         .B(\next_i2c_device_driver_return_state[3] ), .C(\next_i2c_device_driver_state[2] ), 
         .D(n52450), .Z(n47107)) /* synthesis lut_function=(A (C)+!A !((C+(D))+!B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i22_4_lut_4_lut_4_lut_4_lut.init = 16'ha0a4;
    PFUMX i40292 (.BLUT(n51196), .ALUT(n51195), .C0(measurement_period_tx_index[0]), 
          .Z(n51197));
    LUT4 i1_2_lut_rep_476 (.A(resetn), .B(resetn_VL53L1X_buffer), .Z(n52412)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_rep_476.init = 16'h2222;
    LUT4 i1_2_lut_3_lut_adj_344 (.A(resetn), .B(resetn_VL53L1X_buffer), 
         .C(\VL53L1X_data_rx_reg[7] [7]), .Z(VL53L1X_data_rx_reg_7__7__N_473)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_3_lut_adj_344.init = 16'h2020;
    LUT4 i1_2_lut_3_lut_adj_345 (.A(resetn), .B(resetn_VL53L1X_buffer), 
         .C(\VL53L1X_data_rx_reg[5] [0]), .Z(VL53L1X_data_rx_reg_5__0__N_612)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_3_lut_adj_345.init = 16'h2020;
    LUT4 i1_2_lut (.A(\next_i2c_device_driver_state[4] ), .B(data_reg[0]), 
         .Z(n22_adj_5303)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 n37158_bdd_2_lut_40295 (.A(data_tx[4]), .B(\next_i2c_device_driver_state[0] ), 
         .Z(n51133)) /* synthesis lut_function=(A (B)) */ ;
    defparam n37158_bdd_2_lut_40295.init = 16'h8888;
    LUT4 i11614_3_lut_4_lut (.A(n52447), .B(n52218), .C(data_rx[7]), .D(n52364), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[47])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(252[13:59])
    defparam i11614_3_lut_4_lut.init = 16'hfd20;
    LUT4 i12363_3_lut_4_lut (.A(n52447), .B(n52218), .C(data_rx[0]), .D(n52343), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[32])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(252[13:59])
    defparam i12363_3_lut_4_lut.init = 16'hfe10;
    LUT4 i39700_2_lut (.A(\i2c_top_debug[3] ), .B(\i2c_top_debug[4] ), .Z(n49677)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(53[22:35])
    defparam i39700_2_lut.init = 16'hdddd;
    LUT4 i25447_3_lut (.A(cal_reg_addr[4]), .B(data_reg[4]), .C(\next_i2c_device_driver_state[0] ), 
         .Z(n36072)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i25447_3_lut.init = 16'hcaca;
    FD1S3IX i2c_state__i4 (.D(next_i2c_state_4__N_386[3]), .CK(sys_clk), 
            .CD(n53891), .Q(\next_i2c_device_driver_state[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam i2c_state__i4.GSR = "ENABLED";
    FD1S3IX i2c_state__i3 (.D(next_i2c_state_4__N_386[2]), .CK(sys_clk), 
            .CD(n53891), .Q(\next_i2c_device_driver_state[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam i2c_state__i3.GSR = "ENABLED";
    CCU2D add_7877_add_1_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n43986), .S0(n1));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_7877_add_1_cout.INIT0 = 16'h0000;
    defparam add_7877_add_1_cout.INIT1 = 16'h0000;
    defparam add_7877_add_1_cout.INJECT1_0 = "NO";
    defparam add_7877_add_1_cout.INJECT1_1 = "NO";
    FD1S3IX i2c_state__i2 (.D(next_i2c_state_4__N_386[1]), .CK(sys_clk), 
            .CD(n53891), .Q(\next_i2c_device_driver_state[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam i2c_state__i2.GSR = "ENABLED";
    LUT4 i12349_3_lut_4_lut (.A(n52447), .B(n52218), .C(data_rx[1]), .D(n52344), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[33])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(252[13:59])
    defparam i12349_3_lut_4_lut.init = 16'hfe10;
    LUT4 i12347_3_lut_4_lut (.A(n52447), .B(n52218), .C(data_rx[2]), .D(n52345), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[34])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(252[13:59])
    defparam i12347_3_lut_4_lut.init = 16'hfe10;
    LUT4 i12343_3_lut_4_lut (.A(n52447), .B(n52218), .C(data_rx[3]), .D(n52346), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[35])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(252[13:59])
    defparam i12343_3_lut_4_lut.init = 16'hfe10;
    LUT4 led_data_out_4__I_0_859_Mux_6_i21_4_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(data_tx[6]), .C(n53892), .D(next_data_tx_7__N_1024[6]), .Z(n21)) /* synthesis lut_function=(A (B+(C))+!A (C (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam led_data_out_4__I_0_859_Mux_6_i21_4_lut_4_lut.init = 16'hf8a8;
    LUT4 i39575_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52334), 
         .Z(VL53L1X_data_rx_reg_1__1__N_720)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39575_3_lut.init = 16'h5757;
    LUT4 i37709_3_lut_4_lut_4_lut (.A(\next_i2c_device_driver_state[2] ), 
         .B(\next_i2c_device_driver_state[0] ), .C(data_reg[0]), .D(n53892), 
         .Z(n48496)) /* synthesis lut_function=(A (B (C+(D)))+!A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i37709_3_lut_4_lut_4_lut.init = 16'hccc4;
    LUT4 i12329_3_lut_4_lut (.A(n52447), .B(n52218), .C(data_rx[4]), .D(n52347), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[36])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(252[13:59])
    defparam i12329_3_lut_4_lut.init = 16'hfe10;
    LUT4 i12325_3_lut_4_lut (.A(n52447), .B(n52218), .C(data_rx[5]), .D(n52348), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[37])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(252[13:59])
    defparam i12325_3_lut_4_lut.init = 16'hfe10;
    LUT4 i12323_3_lut_4_lut (.A(n52447), .B(n52218), .C(data_rx[6]), .D(n52350), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[38])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(252[13:59])
    defparam i12323_3_lut_4_lut.init = 16'hfe10;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(\next_i2c_device_driver_state[2] ), 
         .B(\next_i2c_device_driver_state[3] ), .C(next_cal_reg_addr_7__N_1124[7]), 
         .D(n52440), .Z(n47981)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'h4000;
    LUT4 i12309_3_lut_4_lut (.A(n52447), .B(n52218), .C(data_rx[7]), .D(n52351), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[39])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(252[13:59])
    defparam i12309_3_lut_4_lut.init = 16'hfe10;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_346 (.A(\next_i2c_device_driver_state[2] ), 
         .B(\next_i2c_device_driver_state[3] ), .C(next_cal_reg_addr_7__N_1124[6]), 
         .D(n52440), .Z(n47983)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_346.init = 16'h4000;
    LUT4 i23_3_lut_3_lut (.A(\next_i2c_device_driver_state[2] ), .B(\next_i2c_device_driver_state[0] ), 
         .C(\next_i2c_device_driver_return_state[3] ), .Z(n9)) /* synthesis lut_function=(A (B (C))+!A ((C)+!B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i23_3_lut_3_lut.init = 16'hd1d1;
    LUT4 i27025_2_lut_4_lut_4_lut (.A(\next_i2c_device_driver_state[2] ), 
         .B(\next_i2c_device_driver_state[3] ), .C(n52177), .D(n3_adj_5304), 
         .Z(n23405)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i27025_2_lut_4_lut_4_lut.init = 16'h5140;
    LUT4 i33204_2_lut (.A(count_ms[0]), .B(count_ms[15]), .Z(n43843)) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i33204_2_lut.init = 16'h9999;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_347 (.A(\next_i2c_device_driver_state[2] ), 
         .B(\next_i2c_device_driver_state[3] ), .C(next_cal_reg_addr_7__N_1124[4]), 
         .D(n52440), .Z(n47982)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_347.init = 16'h4000;
    LUT4 i4_4_lut_rep_534 (.A(n7_adj_5271), .B(n7250), .C(\next_i2c_device_driver_state[0] ), 
         .D(n52210), .Z(n53888)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i4_4_lut_rep_534.init = 16'h8000;
    LUT4 i39827_3_lut (.A(cal_reg_addr[7]), .B(cal_reg_addr[6]), .C(cal_reg_addr[5]), 
         .Z(n49535)) /* synthesis lut_function=(A+!(B (C))) */ ;
    defparam i39827_3_lut.init = 16'hbfbf;
    LUT4 i39464_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52386), 
         .Z(VL53L1X_data_rx_reg_7__6__N_482)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39464_3_lut.init = 16'h5757;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_adj_348 (.A(\next_i2c_device_driver_state[2] ), 
         .B(\next_i2c_device_driver_state[3] ), .C(next_cal_reg_addr_7__N_1124[1]), 
         .D(n52440), .Z(n47980)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i1_2_lut_3_lut_4_lut_4_lut_adj_348.init = 16'h4000;
    LUT4 i2_2_lut_2_lut (.A(\next_i2c_device_driver_state[2] ), .B(n53892), 
         .Z(n7_adj_5301)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i2_2_lut_2_lut.init = 16'h4444;
    LUT4 i12461_3_lut_4_lut (.A(n52447), .B(n52219), .C(data_rx[0]), .D(n52333), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[8])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(229[14] 230[75])
    defparam i12461_3_lut_4_lut.init = 16'hfd20;
    LUT4 i12455_3_lut_4_lut (.A(n52447), .B(n52219), .C(data_rx[1]), .D(n52334), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[9])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(229[14] 230[75])
    defparam i12455_3_lut_4_lut.init = 16'hfd20;
    LUT4 i39467_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52384), 
         .Z(VL53L1X_data_rx_reg_7__5__N_488)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39467_3_lut.init = 16'h5757;
    FD1P3IX master_trigger_count_ms_i5 (.D(n611[5]), .SP(sys_clk_enable_224), 
            .CD(n52182), .CK(sys_clk), .Q(master_trigger_count_ms[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(268[14] 281[12])
    defparam master_trigger_count_ms_i5.GSR = "ENABLED";
    LUT4 i19835_3_lut_rep_393 (.A(n30506), .B(n30505), .C(n30504), .Z(n52329)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19835_3_lut_rep_393.init = 16'hcaca;
    LUT4 i12453_3_lut_4_lut (.A(n52447), .B(n52219), .C(data_rx[2]), .D(n52335), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[10])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(229[14] 230[75])
    defparam i12453_3_lut_4_lut.init = 16'hfd20;
    CCU2D add_7877_add_1_16 (.A0(VL53L1X_osc_cal_val[14]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(VL53L1X_osc_cal_val[15]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n43985), .COUT(n43986), .S0(n2[20]), 
          .S1(n2[21]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_7877_add_1_16.INIT0 = 16'h5aaa;
    defparam add_7877_add_1_16.INIT1 = 16'h5aaa;
    defparam add_7877_add_1_16.INJECT1_0 = "NO";
    defparam add_7877_add_1_16.INJECT1_1 = "NO";
    LUT4 i12449_3_lut_4_lut (.A(n52447), .B(n52219), .C(data_rx[3]), .D(n52336), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[11])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(229[14] 230[75])
    defparam i12449_3_lut_4_lut.init = 16'hfd20;
    FD1P3IX master_trigger_count_ms_i4 (.D(n611[4]), .SP(sys_clk_enable_224), 
            .CD(n52182), .CK(sys_clk), .Q(master_trigger_count_ms[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(268[14] 281[12])
    defparam master_trigger_count_ms_i4.GSR = "ENABLED";
    LUT4 i12439_3_lut_4_lut (.A(n52447), .B(n52219), .C(data_rx[4]), .D(n52337), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[12])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(229[14] 230[75])
    defparam i12439_3_lut_4_lut.init = 16'hfd20;
    CCU2D add_7877_add_1_14 (.A0(VL53L1X_osc_cal_val[12]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(VL53L1X_osc_cal_val[13]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n43984), .COUT(n43985), .S0(n2[18]), 
          .S1(n2[19]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_7877_add_1_14.INIT0 = 16'h5aaa;
    defparam add_7877_add_1_14.INIT1 = 16'h5aaa;
    defparam add_7877_add_1_14.INJECT1_0 = "NO";
    defparam add_7877_add_1_14.INJECT1_1 = "NO";
    CCU2D add_7877_add_1_12 (.A0(VL53L1X_osc_cal_val[10]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(VL53L1X_osc_cal_val[11]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n43983), .COUT(n43984), .S0(n2[16]), 
          .S1(n2[17]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_7877_add_1_12.INIT0 = 16'h5aaa;
    defparam add_7877_add_1_12.INIT1 = 16'h5aaa;
    defparam add_7877_add_1_12.INJECT1_0 = "NO";
    defparam add_7877_add_1_12.INJECT1_1 = "NO";
    LUT4 i39694_2_lut (.A(\next_i2c_device_driver_state[4] ), .B(\next_i2c_device_driver_state[3] ), 
         .Z(n49693)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i39694_2_lut.init = 16'hdddd;
    LUT4 i39470_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52381), 
         .Z(VL53L1X_data_rx_reg_7__4__N_494)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39470_3_lut.init = 16'h5757;
    CCU2D add_7877_add_1_10 (.A0(VL53L1X_osc_cal_val[8]), .B0(VL53L1X_osc_cal_val[14]), 
          .C0(GND_net), .D0(GND_net), .A1(VL53L1X_osc_cal_val[9]), .B1(VL53L1X_osc_cal_val[15]), 
          .C1(GND_net), .D1(GND_net), .CIN(n43982), .COUT(n43983), .S0(n2[14]), 
          .S1(n2[15]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_7877_add_1_10.INIT0 = 16'h5666;
    defparam add_7877_add_1_10.INIT1 = 16'h5666;
    defparam add_7877_add_1_10.INJECT1_0 = "NO";
    defparam add_7877_add_1_10.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut_adj_349 (.A(n30506), .B(n30505), .C(n30504), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_0__4__N_748)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_349.init = 16'hca00;
    LUT4 i11378_3_lut (.A(n52374), .B(data_rx[0]), .C(n28247), .Z(VL53L1X_data_rx_reg_7__7__N_472[56])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i11378_3_lut.init = 16'hcaca;
    LUT4 i19831_3_lut_rep_394 (.A(n30502), .B(n30501), .C(n30500), .Z(n52330)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19831_3_lut_rep_394.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_350 (.A(n30502), .B(n30501), .C(n30500), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_0__5__N_742)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_350.init = 16'hca00;
    LUT4 count_ms_15__I_0_875_i3_3_lut (.A(count_ms_15__N_910[4]), .B(count_ms_15__N_894[2]), 
         .C(n7654[7]), .Z(count_ms_15__N_396[2])) /* synthesis lut_function=(A (B (C))+!A (B+!(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(194[14] 219[12])
    defparam count_ms_15__I_0_875_i3_3_lut.init = 16'hc5c5;
    LUT4 i19827_3_lut_rep_395 (.A(n30498), .B(n30497), .C(n30496), .Z(n52331)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19827_3_lut_rep_395.init = 16'hcaca;
    LUT4 i39473_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52380), 
         .Z(VL53L1X_data_rx_reg_7__3__N_500)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39473_3_lut.init = 16'h5757;
    LUT4 i39448_2_lut_3_lut_4_lut (.A(resetn), .B(wd_event_active), .C(n52515), 
         .D(resetn_imu_N_1182), .Z(sys_clk_enable_256)) /* synthesis lut_function=((B+!(C (D)))+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(371[14:35])
    defparam i39448_2_lut_3_lut_4_lut.init = 16'hdfff;
    FD1P3IX count_ms_i15 (.D(n44[15]), .SP(count_sys_clk_for_ms[16]), .CD(n52172), 
            .CK(sys_clk_N_413), .Q(count_ms[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam count_ms_i15.GSR = "ENABLED";
    FD1P3IX count_ms_i14 (.D(n44[14]), .SP(count_sys_clk_for_ms[16]), .CD(n52172), 
            .CK(sys_clk_N_413), .Q(count_ms[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam count_ms_i14.GSR = "ENABLED";
    FD1P3IX count_ms_i13 (.D(n44[13]), .SP(count_sys_clk_for_ms[16]), .CD(n52172), 
            .CK(sys_clk_N_413), .Q(count_ms[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam count_ms_i13.GSR = "ENABLED";
    FD1P3IX count_ms_i12 (.D(n44[12]), .SP(count_sys_clk_for_ms[16]), .CD(n52172), 
            .CK(sys_clk_N_413), .Q(count_ms[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam count_ms_i12.GSR = "ENABLED";
    FD1P3IX count_ms_i11 (.D(n44[11]), .SP(count_sys_clk_for_ms[16]), .CD(n52172), 
            .CK(sys_clk_N_413), .Q(count_ms[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam count_ms_i11.GSR = "ENABLED";
    FD1P3IX count_ms_i10 (.D(n44[10]), .SP(count_sys_clk_for_ms[16]), .CD(n52172), 
            .CK(sys_clk_N_413), .Q(count_ms[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam count_ms_i10.GSR = "ENABLED";
    FD1P3AY count_ms_i9 (.D(count_ms_15__N_396[9]), .SP(sys_clk_N_413_enable_8), 
            .CK(sys_clk_N_413), .Q(count_ms[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam count_ms_i9.GSR = "ENABLED";
    FD1P3AY count_ms_i8 (.D(count_ms_15__N_396[8]), .SP(sys_clk_N_413_enable_8), 
            .CK(sys_clk_N_413), .Q(count_ms[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam count_ms_i8.GSR = "ENABLED";
    FD1P3AY count_ms_i7 (.D(count_ms_15__N_396[7]), .SP(sys_clk_N_413_enable_8), 
            .CK(sys_clk_N_413), .Q(count_ms[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam count_ms_i7.GSR = "ENABLED";
    LUT4 i39476_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52377), 
         .Z(VL53L1X_data_rx_reg_7__2__N_506)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39476_3_lut.init = 16'h5757;
    LUT4 i1_2_lut_4_lut_adj_351 (.A(n30498), .B(n30497), .C(n30496), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_0__6__N_736)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_351.init = 16'hca00;
    FD1P3AY count_ms_i6 (.D(count_ms_15__N_396[6]), .SP(sys_clk_N_413_enable_8), 
            .CK(sys_clk_N_413), .Q(count_ms[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam count_ms_i6.GSR = "ENABLED";
    FD1P3AY count_ms_i5 (.D(count_ms_15__N_396[5]), .SP(sys_clk_N_413_enable_8), 
            .CK(sys_clk_N_413), .Q(count_ms[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam count_ms_i5.GSR = "ENABLED";
    FD1P3AX count_ms_i4 (.D(count_ms_15__N_396[4]), .SP(sys_clk_N_413_enable_8), 
            .CK(sys_clk_N_413), .Q(count_ms[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam count_ms_i4.GSR = "ENABLED";
    FD1S3AY count_ms_i3 (.D(count_ms_15__N_396[3]), .CK(sys_clk_N_413), 
            .Q(count_ms[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam count_ms_i3.GSR = "ENABLED";
    LUT4 i23_2_lut_rep_484 (.A(\next_i2c_device_driver_state[0] ), .B(n53892), 
         .Z(n52420)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i23_2_lut_rep_484.init = 16'h6666;
    FD1P3AX count_ms_i2 (.D(count_ms_15__N_396[2]), .SP(sys_clk_N_413_enable_8), 
            .CK(sys_clk_N_413), .Q(count_ms[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam count_ms_i2.GSR = "ENABLED";
    LUT4 i26851_2_lut_3_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n53892), .C(data_reg[3]), .D(\next_i2c_device_driver_state[2] ), 
         .Z(n29_adj_5259)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(B (C (D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i26851_2_lut_3_lut_4_lut.init = 16'h6000;
    FD1P3AX count_ms_i1 (.D(count_ms_15__N_396[1]), .SP(sys_clk_N_413_enable_8), 
            .CK(sys_clk_N_413), .Q(count_ms[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam count_ms_i1.GSR = "ENABLED";
    CCU2D add_7877_add_1_8 (.A0(VL53L1X_osc_cal_val[6]), .B0(VL53L1X_osc_cal_val[12]), 
          .C0(GND_net), .D0(GND_net), .A1(VL53L1X_osc_cal_val[7]), .B1(VL53L1X_osc_cal_val[13]), 
          .C1(GND_net), .D1(GND_net), .CIN(n43981), .COUT(n43982), .S0(n2[12]), 
          .S1(n2[13]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_7877_add_1_8.INIT0 = 16'h5666;
    defparam add_7877_add_1_8.INIT1 = 16'h5666;
    defparam add_7877_add_1_8.INJECT1_0 = "NO";
    defparam add_7877_add_1_8.INJECT1_1 = "NO";
    LUT4 i19823_3_lut_rep_396 (.A(n30494), .B(n30493), .C(n30492), .Z(n52332)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19823_3_lut_rep_396.init = 16'hcaca;
    LUT4 i38935_4_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), .B(n53892), 
         .C(\next_i2c_device_driver_state[2] ), .D(data_reg[2]), .Z(n49730)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)))+!A !(B ((D)+!C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i38935_4_lut_4_lut.init = 16'h6c0c;
    LUT4 i1_2_lut_4_lut_adj_352 (.A(n30494), .B(n30493), .C(n30492), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_0__7__N_730)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_352.init = 16'hca00;
    LUT4 i19819_3_lut_rep_397 (.A(n30490), .B(n30489), .C(n30488), .Z(n52333)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19819_3_lut_rep_397.init = 16'hcaca;
    LUT4 i39252_3_lut_3_lut (.A(\next_i2c_device_driver_state[3] ), .B(n52042), 
         .C(n18_adj_5312), .Z(n6_adj_5313)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i39252_3_lut_3_lut.init = 16'he4e4;
    LUT4 i1_2_lut_4_lut_adj_353 (.A(n30490), .B(n30489), .C(n30488), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_1__0__N_724)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_353.init = 16'hca00;
    LUT4 i27012_2_lut_3_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n53892), .C(data_tx[1]), .D(\next_i2c_device_driver_state[2] ), 
         .Z(n29_adj_5266)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(B (C (D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i27012_2_lut_3_lut_4_lut.init = 16'h6000;
    LUT4 i19815_3_lut_rep_398 (.A(n30486), .B(n30485), .C(n30484), .Z(n52334)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19815_3_lut_rep_398.init = 16'hcaca;
    LUT4 i39479_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52376), 
         .Z(VL53L1X_data_rx_reg_7__1__N_512)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39479_3_lut.init = 16'h5757;
    LUT4 i1_2_lut_4_lut_adj_354 (.A(n30486), .B(n30485), .C(n30484), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_1__1__N_718)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_354.init = 16'hca00;
    CCU2D add_409_9 (.A0(cal_reg_addr[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n43786), .S0(next_cal_reg_addr_7__N_1124[7]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(602[42:66])
    defparam add_409_9.INIT0 = 16'h5aaa;
    defparam add_409_9.INIT1 = 16'h0000;
    defparam add_409_9.INJECT1_0 = "NO";
    defparam add_409_9.INJECT1_1 = "NO";
    FD1S3IX data_reg__i8 (.D(next_data_reg_15__N_362[8]), .CK(sys_clk), 
            .CD(n53891), .Q(data_reg[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam data_reg__i8.GSR = "ENABLED";
    LUT4 i1_3_lut (.A(n53892), .B(\next_i2c_device_driver_state[0] ), .C(\next_i2c_state_4__N_1055[1] ), 
         .Z(n33834)) /* synthesis lut_function=(!((B (C))+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam i1_3_lut.init = 16'h2a2a;
    CCU2D add_409_7 (.A0(cal_reg_addr[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cal_reg_addr[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43785), .COUT(n43786), .S0(next_cal_reg_addr_7__N_1124[5]), 
          .S1(next_cal_reg_addr_7__N_1124[6]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(602[42:66])
    defparam add_409_7.INIT0 = 16'h5aaa;
    defparam add_409_7.INIT1 = 16'h5aaa;
    defparam add_409_7.INJECT1_0 = "NO";
    defparam add_409_7.INJECT1_1 = "NO";
    LUT4 i12426_3_lut_4_lut (.A(n52447), .B(n52219), .C(data_rx[5]), .D(n52338), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[13])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(229[14] 230[75])
    defparam i12426_3_lut_4_lut.init = 16'hfd20;
    LUT4 i27146_4_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), .B(n53892), 
         .C(\next_i2c_device_driver_state[2] ), .D(target_read_count[1]), 
         .Z(n14_adj_5314)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C (D))+!B !(C+!(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i27146_4_lut_4_lut.init = 16'h6300;
    LUT4 i19811_3_lut_rep_399 (.A(n30482), .B(n30481), .C(n30480), .Z(n52335)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19811_3_lut_rep_399.init = 16'hcaca;
    LUT4 i13753_2_lut_rep_346_3_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n53892), .C(\next_i2c_device_driver_state[2] ), .Z(n52282)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i13753_2_lut_rep_346_3_lut.init = 16'h6060;
    LUT4 led_data_out_4__I_0_858_Mux_1_i29_4_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n53892), .C(data_reg[1]), .D(\next_i2c_device_driver_state[2] ), 
         .Z(n29_adj_5260)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)))+!A !(B (C+!(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam led_data_out_4__I_0_858_Mux_1_i29_4_lut_4_lut.init = 16'h60cc;
    LUT4 i39482_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52374), 
         .Z(VL53L1X_data_rx_reg_7__0__N_518)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39482_3_lut.init = 16'h5757;
    LUT4 i1_2_lut_4_lut_adj_355 (.A(n30482), .B(n30481), .C(n30480), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_1__2__N_712)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_355.init = 16'hca00;
    LUT4 i19807_3_lut_rep_400 (.A(n30478), .B(n30477), .C(n30476), .Z(n52336)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19807_3_lut_rep_400.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_356 (.A(n30478), .B(n30477), .C(n30476), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_1__3__N_706)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_356.init = 16'hca00;
    FD1S3IX data_reg__i7 (.D(next_data_reg_15__N_362[7]), .CK(sys_clk), 
            .CD(n53891), .Q(data_reg[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam data_reg__i7.GSR = "ENABLED";
    FD1S3IX data_reg__i6 (.D(next_data_reg_15__N_362[6]), .CK(sys_clk), 
            .CD(n53891), .Q(data_reg[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam data_reg__i6.GSR = "ENABLED";
    FD1S3IX data_reg__i5 (.D(next_data_reg_15__N_362[5]), .CK(sys_clk), 
            .CD(n53891), .Q(data_reg[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam data_reg__i5.GSR = "ENABLED";
    CCU2D add_7877_add_1_6 (.A0(VL53L1X_osc_cal_val[4]), .B0(VL53L1X_osc_cal_val[10]), 
          .C0(GND_net), .D0(GND_net), .A1(VL53L1X_osc_cal_val[5]), .B1(VL53L1X_osc_cal_val[11]), 
          .C1(GND_net), .D1(GND_net), .CIN(n43980), .COUT(n43981), .S0(n2[10]), 
          .S1(n2[11]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_7877_add_1_6.INIT0 = 16'h5666;
    defparam add_7877_add_1_6.INIT1 = 16'h5666;
    defparam add_7877_add_1_6.INJECT1_0 = "NO";
    defparam add_7877_add_1_6.INJECT1_1 = "NO";
    CCU2D add_7877_add_1_4 (.A0(VL53L1X_osc_cal_val[2]), .B0(VL53L1X_osc_cal_val[8]), 
          .C0(GND_net), .D0(GND_net), .A1(VL53L1X_osc_cal_val[3]), .B1(VL53L1X_osc_cal_val[9]), 
          .C1(GND_net), .D1(GND_net), .CIN(n43979), .COUT(n43980), .S0(n2[8]), 
          .S1(n2[9]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_7877_add_1_4.INIT0 = 16'h5666;
    defparam add_7877_add_1_4.INIT1 = 16'h5666;
    defparam add_7877_add_1_4.INJECT1_0 = "NO";
    defparam add_7877_add_1_4.INJECT1_1 = "NO";
    CCU2D add_7877_add_1_2 (.A0(VL53L1X_osc_cal_val[0]), .B0(VL53L1X_osc_cal_val[6]), 
          .C0(GND_net), .D0(GND_net), .A1(VL53L1X_osc_cal_val[1]), .B1(VL53L1X_osc_cal_val[7]), 
          .C1(GND_net), .D1(GND_net), .COUT(n43979), .S1(n2[7]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_7877_add_1_2.INIT0 = 16'h7000;
    defparam add_7877_add_1_2.INIT1 = 16'h5666;
    defparam add_7877_add_1_2.INJECT1_0 = "NO";
    defparam add_7877_add_1_2.INJECT1_1 = "NO";
    LUT4 n52078_bdd_4_lut_41628 (.A(n52078), .B(n37158), .C(n19_adj_5319), 
         .D(n53892), .Z(n52134)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A !((D)+!C)) */ ;
    defparam n52078_bdd_4_lut_41628.init = 16'h88f0;
    LUT4 i39938_2_lut_rep_247 (.A(master_trigger_count_ms[20]), .B(n53888), 
         .Z(sys_clk_enable_224)) /* synthesis lut_function=(!(A (B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(273[18:78])
    defparam i39938_2_lut_rep_247.init = 16'h7777;
    LUT4 i1_3_lut_3_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), .B(n53892), 
         .C(data_reg[4]), .D(\next_i2c_device_driver_state[2] ), .Z(n18_adj_5312)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A !(B (C+!(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i1_3_lut_3_lut_4_lut.init = 16'h6066;
    LUT4 i26529_2_lut_3_lut (.A(\next_i2c_device_driver_state[0] ), .B(n53892), 
         .C(data_tx[4]), .Z(n28_adj_5292)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i26529_2_lut_3_lut.init = 16'h6060;
    FD1S3IX data_reg__i4 (.D(next_data_reg_15__N_362[4]), .CK(sys_clk), 
            .CD(n52212), .Q(data_reg[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam data_reg__i4.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_adj_357 (.A(\next_i2c_device_driver_state[0] ), .B(n53892), 
         .C(data_tx[3]), .Z(n19_adj_5281)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i1_2_lut_3_lut_adj_357.init = 16'h6060;
    FD1S3IX data_reg__i3 (.D(next_data_reg_15__N_362[3]), .CK(sys_clk), 
            .CD(n52212), .Q(data_reg[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam data_reg__i3.GSR = "ENABLED";
    FD1S3IX data_reg__i2 (.D(next_data_reg_15__N_362[2]), .CK(sys_clk), 
            .CD(n52212), .Q(data_reg[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam data_reg__i2.GSR = "ENABLED";
    FD1S3IX data_reg__i1 (.D(next_data_reg_15__N_362[1]), .CK(sys_clk), 
            .CD(n52212), .Q(data_reg[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam data_reg__i1.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_adj_358 (.A(\next_i2c_device_driver_state[0] ), .B(n53892), 
         .C(data_tx[7]), .Z(n19_adj_5284)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i1_2_lut_3_lut_adj_358.init = 16'h6060;
    LUT4 i19803_3_lut_rep_401 (.A(n30474), .B(n30473), .C(n30472), .Z(n52337)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19803_3_lut_rep_401.init = 16'hcaca;
    LUT4 i12424_3_lut_4_lut (.A(n52447), .B(n52219), .C(data_rx[6]), .D(n52339), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[14])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(229[14] 230[75])
    defparam i12424_3_lut_4_lut.init = 16'hfd20;
    PFUMX i40247 (.BLUT(n51130), .ALUT(n51129), .C0(measurement_period_tx_index[0]), 
          .Z(n51131));
    LUT4 i1_2_lut_4_lut_adj_359 (.A(n30474), .B(n30473), .C(n30472), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_1__4__N_700)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_359.init = 16'hca00;
    LUT4 i19799_3_lut_rep_402 (.A(n30470), .B(n30469), .C(n30468), .Z(n52338)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19799_3_lut_rep_402.init = 16'hcaca;
    LUT4 i25645_2_lut_3_lut (.A(\next_i2c_device_driver_state[0] ), .B(n53892), 
         .C(data_tx[5]), .Z(n28)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i25645_2_lut_3_lut.init = 16'h6060;
    LUT4 i39485_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52372), 
         .Z(VL53L1X_data_rx_reg_6__7__N_524)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39485_3_lut.init = 16'h5757;
    LUT4 i18385_1_lut_rep_236 (.A(n7654[7]), .Z(n52172)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam i18385_1_lut_rep_236.init = 16'h5555;
    LUT4 i11_4_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), .B(n53892), 
         .C(data_reg[0]), .D(\next_i2c_device_driver_state[4] ), .Z(n46521)) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)))+!A !(B (C+!(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i11_4_lut_4_lut.init = 16'h60cc;
    LUT4 VL53L1X_measurement_period_1__bdd_2_lut_40448 (.A(VL53L1X_measurement_period[9]), 
         .B(measurement_period_tx_index[1]), .Z(n51195)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam VL53L1X_measurement_period_1__bdd_2_lut_40448.init = 16'h2222;
    LUT4 i39488_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52371), 
         .Z(VL53L1X_data_rx_reg_6__6__N_530)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39488_3_lut.init = 16'h5757;
    LUT4 i1_2_lut_4_lut_adj_360 (.A(n30470), .B(n30469), .C(n30468), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_1__5__N_694)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_360.init = 16'hca00;
    LUT4 i2_4_lut (.A(\next_i2c_device_driver_state[2] ), .B(\next_i2c_device_driver_state[0] ), 
         .C(n53892), .D(\next_i2c_device_driver_return_state[3] ), .Z(n48658)) /* synthesis lut_function=(A (B (C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam i2_4_lut.init = 16'h8880;
    LUT4 i19795_3_lut_rep_403 (.A(n30466), .B(n30465), .C(n30464), .Z(n52339)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19795_3_lut_rep_403.init = 16'hcaca;
    FD1P3IX master_trigger_count_ms_i3 (.D(n611[3]), .SP(sys_clk_enable_224), 
            .CD(n52182), .CK(sys_clk), .Q(master_trigger_count_ms[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(268[14] 281[12])
    defparam master_trigger_count_ms_i3.GSR = "ENABLED";
    LUT4 mux_833_Mux_4_i127_4_lut (.A(n28179), .B(n47344), .C(cal_reg_addr[7]), 
         .D(n47394), .Z(n127)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (B+!(C)))) */ ;
    defparam mux_833_Mux_4_i127_4_lut.init = 16'h3a30;
    LUT4 i17669_2_lut (.A(cal_reg_addr[0]), .B(cal_reg_addr[3]), .Z(n28179)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i17669_2_lut.init = 16'h6666;
    LUT4 i38928_4_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), .B(n53892), 
         .C(\next_i2c_device_driver_state[2] ), .D(data_reg[7]), .Z(n49723)) /* synthesis lut_function=(!(A (B (C)+!B !(C (D)))+!A !(B ((D)+!C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i38928_4_lut_4_lut.init = 16'h6c0c;
    LUT4 i26045_2_lut_3_lut (.A(\next_i2c_device_driver_state[0] ), .B(n53892), 
         .C(data_tx[2]), .Z(n28_adj_5279)) /* synthesis lut_function=(!(A (B+!(C))+!A !(B (C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i26045_2_lut_3_lut.init = 16'h6060;
    LUT4 i24317_1_lut_rep_485 (.A(\next_i2c_device_driver_state[0] ), .Z(n52421)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam i24317_1_lut_rep_485.init = 16'h5555;
    LUT4 i1_2_lut_3_lut_4_lut_4_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n53892), .C(n53056), .D(\next_i2c_device_driver_state[2] ), 
         .Z(n30_adj_5320)) /* synthesis lut_function=(A (C)+!A (B (C+!(D))+!B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam i1_2_lut_3_lut_4_lut_4_lut_4_lut.init = 16'hf0f4;
    LUT4 i39491_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52370), 
         .Z(VL53L1X_data_rx_reg_6__5__N_536)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39491_3_lut.init = 16'h5757;
    LUT4 i23188_3_lut_4_lut_4_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(\next_i2c_device_driver_return_state[0] ), .C(\next_i2c_device_driver_state[4] ), 
         .D(n52283), .Z(n33840)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C+!(D))+!B (C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam i23188_3_lut_4_lut_4_lut_4_lut.init = 16'h505c;
    LUT4 i12422_3_lut_4_lut (.A(n52447), .B(n52219), .C(data_rx[7]), .D(n52340), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[15])) /* synthesis lut_function=(A (B (D)+!B (C))+!A (D)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(229[14] 230[75])
    defparam i12422_3_lut_4_lut.init = 16'hfd20;
    LUT4 i2_4_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), .B(n21_adj_5321), 
         .C(n49547), .D(n24_adj_5322), .Z(n7246)) /* synthesis lut_function=(A (B+(D))+!A (B+((D)+!C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam i2_4_lut_4_lut.init = 16'hffcd;
    LUT4 i11371_3_lut (.A(n52376), .B(data_rx[1]), .C(n28247), .Z(VL53L1X_data_rx_reg_7__7__N_472[57])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i11371_3_lut.init = 16'hcaca;
    CCU2D add_8435_22 (.A0(n2[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n1), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n43976), 
          .S0(n25[21]), .S1(n25[22]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_8435_22.INIT0 = 16'h5aaa;
    defparam add_8435_22.INIT1 = 16'h5aaa;
    defparam add_8435_22.INJECT1_0 = "NO";
    defparam add_8435_22.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut_adj_361 (.A(n30466), .B(n30465), .C(n30464), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_1__6__N_688)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_361.init = 16'hca00;
    LUT4 i1_3_lut_4_lut_3_lut (.A(\next_i2c_device_driver_state[0] ), .B(cal_reg_addr[5]), 
         .C(data_reg[5]), .Z(n8_adj_5323)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam i1_3_lut_4_lut_3_lut.init = 16'he4e4;
    LUT4 i26146_4_lut_4_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n1_adj_5324), .C(n53892), .D(\next_i2c_device_driver_state[2] ), 
         .Z(n7_adj_5325)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (B (D)+!B ((D)+!C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam i26146_4_lut_4_lut_4_lut.init = 16'h005c;
    LUT4 VL53L1X_measurement_period_1__bdd_3_lut_40449 (.A(VL53L1X_measurement_period[1]), 
         .B(measurement_period_tx_index[1]), .C(VL53L1X_measurement_period[17]), 
         .Z(n51196)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam VL53L1X_measurement_period_1__bdd_3_lut_40449.init = 16'he2e2;
    LUT4 i19791_3_lut_rep_404 (.A(n30462), .B(n30461), .C(n30460), .Z(n52340)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19791_3_lut_rep_404.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_362 (.A(n30462), .B(n30461), .C(n30460), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_1__7__N_682)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_362.init = 16'hca00;
    LUT4 i39494_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52369), 
         .Z(VL53L1X_data_rx_reg_6__4__N_542)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39494_3_lut.init = 16'h5757;
    LUT4 i11158_3_lut_4_lut (.A(n52447), .B(n52219), .C(data_rx[0]), .D(n52320), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[0])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(229[14] 230[75])
    defparam i11158_3_lut_4_lut.init = 16'hfe10;
    LUT4 i39328_4_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), .B(n49637), 
         .C(next_data_tx_7__N_1032_c[4]), .D(n126), .Z(n8_adj_5326)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam i39328_4_lut_4_lut.init = 16'hf4b0;
    LUT4 i10_then_4_lut (.A(\next_i2c_device_driver_state[3] ), .B(n53892), 
         .C(\next_i2c_device_driver_state[4] ), .D(\next_i2c_device_driver_state[2] ), 
         .Z(n52499)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (C+!(D)))) */ ;
    defparam i10_then_4_lut.init = 16'h0508;
    LUT4 n37158_bdd_2_lut_40326 (.A(data_tx[1]), .B(\next_i2c_device_driver_state[0] ), 
         .Z(n51199)) /* synthesis lut_function=(A (B)) */ ;
    defparam n37158_bdd_2_lut_40326.init = 16'h8888;
    LUT4 n14_bdd_3_lut_4_lut_4_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n53892), .C(data_reg[4]), .D(\next_i2c_device_driver_state[2] ), 
         .Z(n52040)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B+!(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam n14_bdd_3_lut_4_lut_4_lut_4_lut.init = 16'h3100;
    LUT4 led_data_out_4__I_0_860_Mux_1_i28_4_lut_3_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n52188), .C(n53892), .Z(n28_adj_5327)) /* synthesis lut_function=(!(A (B+(C))+!A !(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam led_data_out_4__I_0_860_Mux_1_i28_4_lut_3_lut.init = 16'h5252;
    LUT4 i11330_3_lut_4_lut (.A(n52447), .B(n52219), .C(data_rx[1]), .D(n52321), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[1])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(229[14] 230[75])
    defparam i11330_3_lut_4_lut.init = 16'hfe10;
    LUT4 i1_3_lut_4_lut_3_lut_adj_363 (.A(\next_i2c_device_driver_state[0] ), 
         .B(next_data_tx_7__N_1032_c[6]), .C(data_tx[6]), .Z(n8)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam i1_3_lut_4_lut_3_lut_adj_363.init = 16'he4e4;
    LUT4 i39497_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52368), 
         .Z(VL53L1X_data_rx_reg_6__3__N_548)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39497_3_lut.init = 16'h5757;
    LUT4 i39500_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52367), 
         .Z(VL53L1X_data_rx_reg_6__2__N_554)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39500_3_lut.init = 16'h5757;
    LUT4 led_data_out_4__I_0_859_Mux_0_i22_4_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n53892), .C(\next_i2c_device_driver_state[2] ), .D(n52134), 
         .Z(n22_adj_5328)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A ((D)+!C)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam led_data_out_4__I_0_859_Mux_0_i22_4_lut_4_lut.init = 16'hfd0d;
    LUT4 i1_2_lut_rep_297_3_lut_3_lut_3_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n53892), .C(\next_i2c_device_driver_state[2] ), .Z(n52233)) /* synthesis lut_function=((B+!(C))+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam i1_2_lut_rep_297_3_lut_3_lut_3_lut.init = 16'hdfdf;
    CCU2D add_8435_20 (.A0(n2[19]), .B0(n17827), .C0(GND_net), .D0(GND_net), 
          .A1(n2[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n43975), 
          .COUT(n43976), .S0(n25[19]), .S1(n25[20]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_8435_20.INIT0 = 16'h5666;
    defparam add_8435_20.INIT1 = 16'h5aaa;
    defparam add_8435_20.INJECT1_0 = "NO";
    defparam add_8435_20.INJECT1_1 = "NO";
    CCU2D add_8435_18 (.A0(n2[17]), .B0(n17807[17]), .C0(GND_net), .D0(GND_net), 
          .A1(n2[18]), .B1(n17807[18]), .C1(GND_net), .D1(GND_net), 
          .CIN(n43974), .COUT(n43975), .S0(n25[17]), .S1(n25[18]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_8435_18.INIT0 = 16'h5666;
    defparam add_8435_18.INIT1 = 16'h5666;
    defparam add_8435_18.INJECT1_0 = "NO";
    defparam add_8435_18.INJECT1_1 = "NO";
    LUT4 i39300_3_lut_4_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n13144[4]), .C(n7246), .D(n7240), .Z(n13181[4])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B+!(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam i39300_3_lut_4_lut_4_lut.init = 16'hcfc5;
    CCU2D add_8435_16 (.A0(n2[15]), .B0(n17807[15]), .C0(GND_net), .D0(GND_net), 
          .A1(n2[16]), .B1(n17807[16]), .C1(GND_net), .D1(GND_net), 
          .CIN(n43973), .COUT(n43974), .S0(n25[15]), .S1(n25[16]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_8435_16.INIT0 = 16'h5666;
    defparam add_8435_16.INIT1 = 16'h5666;
    defparam add_8435_16.INJECT1_0 = "NO";
    defparam add_8435_16.INJECT1_1 = "NO";
    LUT4 i1_4_lut_4_lut_adj_364 (.A(\next_i2c_device_driver_state[0] ), .B(n24_adj_5322), 
         .C(n7240), .D(n21_adj_5321), .Z(n48822)) /* synthesis lut_function=((B+(C+(D)))+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam i1_4_lut_4_lut_adj_364.init = 16'hfffd;
    LUT4 i39503_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52366), 
         .Z(VL53L1X_data_rx_reg_6__1__N_560)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39503_3_lut.init = 16'h5757;
    LUT4 i1_4_lut_4_lut_adj_365 (.A(\next_i2c_device_driver_state[0] ), .B(n52460), 
         .C(n7_adj_5301), .D(n53890), .Z(n6974)) /* synthesis lut_function=(A (D)+!A (B (C+(D))+!B (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam i1_4_lut_4_lut_adj_365.init = 16'hff40;
    LUT4 i11280_3_lut_4_lut (.A(n52447), .B(n52219), .C(data_rx[2]), .D(n52322), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[2])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(229[14] 230[75])
    defparam i11280_3_lut_4_lut.init = 16'hfe10;
    LUT4 i20055_2_lut_3_lut_2_lut (.A(master_trigger_count_ms[20]), .B(n53888), 
         .Z(n52182)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(273[18:78])
    defparam i20055_2_lut_3_lut_2_lut.init = 16'h2222;
    LUT4 i13888_4_lut_4_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(data_reg[1]), .C(n53892), .D(\next_i2c_device_driver_state[2] ), 
         .Z(n24343)) /* synthesis lut_function=(A (B+(C+!(D)))+!A !(C)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam i13888_4_lut_4_lut_4_lut.init = 16'hadaf;
    LUT4 mux_833_Mux_4_i255_3_lut (.A(n127), .B(data_tx[4]), .C(\next_i2c_device_driver_state[0] ), 
         .Z(next_data_tx_7__N_1032_c[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam mux_833_Mux_4_i255_3_lut.init = 16'hcaca;
    LUT4 i39506_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52365), 
         .Z(VL53L1X_data_rx_reg_6__0__N_566)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39506_3_lut.init = 16'h5757;
    LUT4 i12943_3_lut_4_lut (.A(n52447), .B(n52219), .C(data_rx[3]), .D(n52324), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[3])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(229[14] 230[75])
    defparam i12943_3_lut_4_lut.init = 16'hfe10;
    LUT4 i12832_3_lut_4_lut (.A(n52447), .B(n52219), .C(data_rx[4]), .D(n52329), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[4])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(229[14] 230[75])
    defparam i12832_3_lut_4_lut.init = 16'hfe10;
    CCU2D add_8435_14 (.A0(n2[13]), .B0(n17807[13]), .C0(GND_net), .D0(GND_net), 
          .A1(n2[14]), .B1(n17807[14]), .C1(GND_net), .D1(GND_net), 
          .CIN(n43972), .COUT(n43973), .S0(n25[13]), .S1(n25[14]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_8435_14.INIT0 = 16'h5666;
    defparam add_8435_14.INIT1 = 16'h5666;
    defparam add_8435_14.INJECT1_0 = "NO";
    defparam add_8435_14.INJECT1_1 = "NO";
    LUT4 i10_else_4_lut (.A(\next_i2c_device_driver_state[3] ), .B(n53892), 
         .C(\next_i2c_device_driver_state[4] ), .D(\next_i2c_device_driver_state[2] ), 
         .Z(n52498)) /* synthesis lut_function=(!(A (B (C+(D))+!B (C (D)+!C !(D)))+!A ((C+!(D))+!B))) */ ;
    defparam i10_else_4_lut.init = 16'h0628;
    CCU2D add_8435_12 (.A0(n2[11]), .B0(n17807[11]), .C0(GND_net), .D0(GND_net), 
          .A1(n2[12]), .B1(n17807[12]), .C1(GND_net), .D1(GND_net), 
          .CIN(n43971), .COUT(n43972), .S0(n25[11]), .S1(n25[12]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_8435_12.INIT0 = 16'h5666;
    defparam add_8435_12.INIT1 = 16'h5666;
    defparam add_8435_12.INJECT1_0 = "NO";
    defparam add_8435_12.INJECT1_1 = "NO";
    LUT4 n53053_bdd_3_lut (.A(n53053), .B(n53050), .C(n53892), .Z(n53054)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n53053_bdd_3_lut.init = 16'hcaca;
    LUT4 next_i2c_device_driver_state_1__bdd_3_lut_41285 (.A(n53892), .B(\next_i2c_device_driver_state[2] ), 
         .C(\next_i2c_device_driver_state[0] ), .Z(n53055)) /* synthesis lut_function=(A+!(B (C))) */ ;
    defparam next_i2c_device_driver_state_1__bdd_3_lut_41285.init = 16'hbfbf;
    LUT4 i19787_3_lut_rep_407 (.A(n30458), .B(n30457), .C(n30456), .Z(n52343)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19787_3_lut_rep_407.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_366 (.A(n30458), .B(n30457), .C(n30456), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_4__0__N_660)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_366.init = 16'hca00;
    LUT4 i1_2_lut_2_lut (.A(n7654[7]), .B(count_sys_clk_for_ms[16]), .Z(sys_clk_N_413_enable_8)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam i1_2_lut_2_lut.init = 16'hdddd;
    LUT4 i25983_4_lut_then_3_lut (.A(cal_reg_addr[4]), .B(cal_reg_addr[1]), 
         .C(cal_reg_addr[0]), .Z(n52502)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i25983_4_lut_then_3_lut.init = 16'h8080;
    LUT4 i38638_4_lut_4_lut (.A(n53892), .B(n33834), .C(\next_i2c_device_driver_state[2] ), 
         .D(n38), .Z(n49433)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (B+((D)+!C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i38638_4_lut_4_lut.init = 16'hf5c5;
    LUT4 i12814_3_lut_4_lut (.A(n52447), .B(n52219), .C(data_rx[5]), .D(n52330), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[5])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(229[14] 230[75])
    defparam i12814_3_lut_4_lut.init = 16'hfe10;
    LUT4 i27175_2_lut_4_lut_4_lut (.A(n53892), .B(\next_i2c_device_driver_state[2] ), 
         .C(n11_adj_5331), .D(n52209), .Z(n22527)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i27175_2_lut_4_lut_4_lut.init = 16'h5140;
    LUT4 i12771_3_lut_4_lut (.A(n52447), .B(n52219), .C(data_rx[6]), .D(n52331), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[6])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(229[14] 230[75])
    defparam i12771_3_lut_4_lut.init = 16'hfe10;
    LUT4 i1_4_lut_4_lut_adj_367 (.A(n53892), .B(\next_i2c_device_driver_state[0] ), 
         .C(n22_adj_5303), .D(n5_adj_5332), .Z(n6_adj_5333)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i1_4_lut_4_lut_adj_367.init = 16'h5140;
    LUT4 i12491_3_lut_4_lut (.A(n52447), .B(n52219), .C(data_rx[7]), .D(n52332), 
         .Z(VL53L1X_data_rx_reg_7__7__N_472[7])) /* synthesis lut_function=(A (D)+!A (B (D)+!B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(229[14] 230[75])
    defparam i12491_3_lut_4_lut.init = 16'hfe10;
    LUT4 i39509_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52364), 
         .Z(VL53L1X_data_rx_reg_5__7__N_572)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39509_3_lut.init = 16'h5757;
    LUT4 i25971_2_lut_2_lut (.A(n7654[7]), .B(count_ms_15__N_894[1]), .Z(count_ms_15__N_396[1])) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam i25971_2_lut_2_lut.init = 16'hdddd;
    LUT4 i19783_3_lut_rep_408 (.A(n30454), .B(n30453), .C(n30452), .Z(n52344)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19783_3_lut_rep_408.init = 16'hcaca;
    LUT4 i39512_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52363), 
         .Z(VL53L1X_data_rx_reg_5__6__N_578)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39512_3_lut.init = 16'h5757;
    LUT4 i26565_2_lut_rep_241_2_lut (.A(n53892), .B(n8_adj_5326), .Z(n52177)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i26565_2_lut_rep_241_2_lut.init = 16'h4444;
    PFUMX i40226 (.BLUT(n51100), .ALUT(n51099), .C0(measurement_period_tx_index[0]), 
          .Z(n51101));
    LUT4 i39836_4_lut (.A(next_addr_7__N_1168), .B(n2485[7]), .C(n52248), 
         .D(n49226), .Z(n48986)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam i39836_4_lut.init = 16'h0020;
    LUT4 i1_2_lut_4_lut_adj_368 (.A(n30454), .B(n30453), .C(n30452), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_4__1__N_654)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_368.init = 16'hca00;
    LUT4 i19779_3_lut_rep_409 (.A(n30450), .B(n30449), .C(n30448), .Z(n52345)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19779_3_lut_rep_409.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_369 (.A(n30450), .B(n30449), .C(n30448), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_4__2__N_648)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_369.init = 16'hca00;
    LUT4 i39515_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52360), 
         .Z(VL53L1X_data_rx_reg_5__5__N_584)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39515_3_lut.init = 16'h5757;
    LUT4 i26145_2_lut_rep_273_4_lut (.A(n52274), .B(cal_reg_addr[7]), .C(n27913), 
         .D(\next_i2c_device_driver_state[0] ), .Z(n52209)) /* synthesis lut_function=(A (B (D))+!A (B (C (D)))) */ ;
    defparam i26145_2_lut_rep_273_4_lut.init = 16'hc800;
    LUT4 i25983_4_lut_else_3_lut (.A(cal_reg_addr[4]), .B(cal_reg_addr[1]), 
         .C(cal_reg_addr[0]), .D(cal_reg_addr[3]), .Z(n52501)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i25983_4_lut_else_3_lut.init = 16'h0200;
    LUT4 i26650_2_lut_3_lut_4_lut (.A(resetn), .B(wd_event_active), .C(n2485[4]), 
         .D(resetn_imu_N_1182), .Z(n7654[4])) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(371[14:35])
    defparam i26650_2_lut_3_lut_4_lut.init = 16'h2000;
    LUT4 i26175_3_lut_3_lut_3_lut (.A(n53892), .B(n52227), .C(\next_i2c_device_driver_state[0] ), 
         .Z(n10_adj_5286)) /* synthesis lut_function=(!(A+!(B+!(C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i26175_3_lut_3_lut_3_lut.init = 16'h4545;
    LUT4 i39518_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52358), 
         .Z(VL53L1X_data_rx_reg_5__4__N_590)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39518_3_lut.init = 16'h5757;
    LUT4 i1_4_lut_4_lut_4_lut_adj_370 (.A(n53892), .B(\next_i2c_device_driver_state[2] ), 
         .C(data_reg[6]), .D(\next_i2c_device_driver_state[0] ), .Z(n47057)) /* synthesis lut_function=(!(A ((D)+!B)+!A !(B (C+!(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i1_4_lut_4_lut_4_lut_adj_370.init = 16'h40cc;
    LUT4 i2_4_lut_4_lut_adj_371 (.A(n53892), .B(\next_i2c_device_driver_state[0] ), 
         .C(measurement_period_tx_index[0]), .D(n53890), .Z(next_measurement_period_tx_index[0])) /* synthesis lut_function=((B (C+(D))+!B ((D)+!C))+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i2_4_lut_4_lut_adj_371.init = 16'hffd7;
    LUT4 i39721_2_lut_rep_295_4_lut_4_lut (.A(n53892), .B(n52303), .C(n52409), 
         .D(n52410), .Z(n52231)) /* synthesis lut_function=(!(A (B)+!A (B+(C (D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i39721_2_lut_rep_295_4_lut_4_lut.init = 16'h2333;
    LUT4 i2_3_lut_rep_344_4_lut_4_lut (.A(n53892), .B(n52410), .C(\next_i2c_device_driver_state[4] ), 
         .D(\next_i2c_device_driver_state[0] ), .Z(sys_clk_enable_108)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i2_3_lut_rep_344_4_lut_4_lut.init = 16'h4000;
    LUT4 i19_4_lut_4_lut_4_lut (.A(n53892), .B(data_reg[3]), .C(\next_i2c_device_driver_state[2] ), 
         .D(\next_i2c_device_driver_state[0] ), .Z(n47071)) /* synthesis lut_function=(!(A (C (D))+!A !(B (C)+!B !((D)+!C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i19_4_lut_4_lut_4_lut.init = 16'h4afa;
    CCU2D add_8435_10 (.A0(n2[9]), .B0(n17807[9]), .C0(GND_net), .D0(GND_net), 
          .A1(n2[10]), .B1(n17807[10]), .C1(GND_net), .D1(GND_net), 
          .CIN(n43970), .COUT(n43971), .S0(n25[9]), .S1(n25[10]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_8435_10.INIT0 = 16'h5666;
    defparam add_8435_10.INIT1 = 16'h5666;
    defparam add_8435_10.INJECT1_0 = "NO";
    defparam add_8435_10.INJECT1_1 = "NO";
    LUT4 i37_then_4_lut (.A(n53892), .B(\next_i2c_device_driver_state[0] ), 
         .C(\next_i2c_device_driver_state[3] ), .D(\next_i2c_device_driver_state[4] ), 
         .Z(n52514)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (B (C+(D))+!B (C (D)))) */ ;
    defparam i37_then_4_lut.init = 16'hfe60;
    CCU2D add_8435_8 (.A0(n2[7]), .B0(n17807[7]), .C0(GND_net), .D0(GND_net), 
          .A1(n2[8]), .B1(n17807[8]), .C1(GND_net), .D1(GND_net), .CIN(n43969), 
          .COUT(n43970), .S0(n25[7]), .S1(n25[8]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_8435_8.INIT0 = 16'h5666;
    defparam add_8435_8.INIT1 = 16'h5666;
    defparam add_8435_8.INJECT1_0 = "NO";
    defparam add_8435_8.INJECT1_1 = "NO";
    CCU2D add_8435_6 (.A0(VL53L1X_osc_cal_val[5]), .B0(n17807[5]), .C0(GND_net), 
          .D0(GND_net), .A1(n2[6]), .B1(n17807[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n43968), .COUT(n43969), .S0(n25[5]), .S1(n25[6]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_8435_6.INIT0 = 16'h5666;
    defparam add_8435_6.INIT1 = 16'h5666;
    defparam add_8435_6.INJECT1_0 = "NO";
    defparam add_8435_6.INJECT1_1 = "NO";
    CCU2D add_8435_4 (.A0(VL53L1X_osc_cal_val[2]), .B0(VL53L1X_osc_cal_val[0]), 
          .C0(VL53L1X_osc_cal_val[3]), .D0(GND_net), .A1(VL53L1X_osc_cal_val[4]), 
          .B1(n17807[4]), .C1(GND_net), .D1(GND_net), .CIN(n43967), 
          .COUT(n43968), .S0(next_VL53L1X_measurement_period_31__N_1103[3]), 
          .S1(next_VL53L1X_measurement_period_31__N_1103[4]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_8435_4.INIT0 = 16'h9696;
    defparam add_8435_4.INIT1 = 16'h5666;
    defparam add_8435_4.INJECT1_0 = "NO";
    defparam add_8435_4.INJECT1_1 = "NO";
    LUT4 i19775_3_lut_rep_410 (.A(n30446), .B(n30445), .C(n30444), .Z(n52346)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19775_3_lut_rep_410.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_372 (.A(n30446), .B(n30445), .C(n30444), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_4__3__N_642)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_372.init = 16'hca00;
    LUT4 i19771_3_lut_rep_411 (.A(n30442), .B(n30441), .C(n30440), .Z(n52347)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19771_3_lut_rep_411.init = 16'hcaca;
    LUT4 i39521_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52357), 
         .Z(VL53L1X_data_rx_reg_5__3__N_596)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39521_3_lut.init = 16'h5757;
    LUT4 i1_2_lut_4_lut_adj_373 (.A(n30442), .B(n30441), .C(n30440), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_4__4__N_636)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_373.init = 16'hca00;
    LUT4 i2_4_lut_then_4_lut (.A(cal_reg_addr[4]), .B(cal_reg_addr[2]), 
         .C(cal_reg_addr[3]), .D(cal_reg_addr[1]), .Z(n52505)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i2_4_lut_then_4_lut.init = 16'h0010;
    LUT4 i19767_3_lut_rep_412 (.A(n30438), .B(n30437), .C(n30436), .Z(n52348)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19767_3_lut_rep_412.init = 16'hcaca;
    FD1P3AX VL53L1X_chip_id_i0_i1 (.D(n52334), .SP(sys_clk_enable_123), 
            .CK(sys_clk), .Q(next_VL53L1X_chip_id[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_chip_id_i0_i1.GSR = "ENABLED";
    FD1P3AX VL53L1X_chip_id_i0_i2 (.D(n52335), .SP(n7654[6]), .CK(sys_clk), 
            .Q(next_VL53L1X_chip_id[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_chip_id_i0_i2.GSR = "ENABLED";
    FD1P3AX VL53L1X_chip_id_i0_i3 (.D(n52336), .SP(n7654[6]), .CK(sys_clk), 
            .Q(next_VL53L1X_chip_id[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_chip_id_i0_i3.GSR = "ENABLED";
    FD1P3AX VL53L1X_chip_id_i0_i4 (.D(n52337), .SP(n7654[6]), .CK(sys_clk), 
            .Q(next_VL53L1X_chip_id[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_chip_id_i0_i4.GSR = "ENABLED";
    FD1P3AX VL53L1X_chip_id_i0_i5 (.D(n52338), .SP(n7654[6]), .CK(sys_clk), 
            .Q(next_VL53L1X_chip_id[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_chip_id_i0_i5.GSR = "ENABLED";
    FD1P3AX VL53L1X_chip_id_i0_i6 (.D(n52339), .SP(n7654[6]), .CK(sys_clk), 
            .Q(next_VL53L1X_chip_id[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_chip_id_i0_i6.GSR = "ENABLED";
    FD1P3AX VL53L1X_chip_id_i0_i7 (.D(n52340), .SP(n7654[6]), .CK(sys_clk), 
            .Q(next_VL53L1X_chip_id[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_chip_id_i0_i7.GSR = "ENABLED";
    FD1P3AX VL53L1X_chip_id_i0_i8 (.D(n52320), .SP(n7654[6]), .CK(sys_clk), 
            .Q(next_VL53L1X_chip_id[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_chip_id_i0_i8.GSR = "ENABLED";
    FD1P3AX VL53L1X_chip_id_i0_i9 (.D(n52321), .SP(n7654[6]), .CK(sys_clk), 
            .Q(next_VL53L1X_chip_id[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_chip_id_i0_i9.GSR = "ENABLED";
    FD1P3AX VL53L1X_chip_id_i0_i10 (.D(n52322), .SP(n7654[6]), .CK(sys_clk), 
            .Q(next_VL53L1X_chip_id[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_chip_id_i0_i10.GSR = "ENABLED";
    FD1P3AX VL53L1X_chip_id_i0_i11 (.D(n52324), .SP(n7654[6]), .CK(sys_clk), 
            .Q(next_VL53L1X_chip_id[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_chip_id_i0_i11.GSR = "ENABLED";
    FD1P3AX VL53L1X_chip_id_i0_i12 (.D(n52329), .SP(n7654[6]), .CK(sys_clk), 
            .Q(next_VL53L1X_chip_id[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_chip_id_i0_i12.GSR = "ENABLED";
    FD1P3AX VL53L1X_chip_id_i0_i13 (.D(n52330), .SP(n7654[6]), .CK(sys_clk), 
            .Q(next_VL53L1X_chip_id[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_chip_id_i0_i13.GSR = "ENABLED";
    FD1P3AX VL53L1X_chip_id_i0_i14 (.D(n52331), .SP(n7654[6]), .CK(sys_clk), 
            .Q(next_VL53L1X_chip_id[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_chip_id_i0_i14.GSR = "ENABLED";
    FD1P3AX VL53L1X_chip_id_i0_i15 (.D(n52332), .SP(n7654[6]), .CK(sys_clk), 
            .Q(next_VL53L1X_chip_id[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(317[14] 323[12])
    defparam VL53L1X_chip_id_i0_i15.GSR = "ENABLED";
    LUT4 i1_2_lut_4_lut_adj_374 (.A(n30438), .B(n30437), .C(n30436), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_4__5__N_630)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_374.init = 16'hca00;
    LUT4 i11369_3_lut (.A(n52377), .B(data_rx[2]), .C(n28247), .Z(VL53L1X_data_rx_reg_7__7__N_472[58])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i11369_3_lut.init = 16'hcaca;
    LUT4 i2_4_lut_else_4_lut (.A(cal_reg_addr[4]), .B(cal_reg_addr[2]), 
         .C(cal_reg_addr[3]), .D(cal_reg_addr[1]), .Z(n52504)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i2_4_lut_else_4_lut.init = 16'h0100;
    LUT4 led_data_out_4__I_0_858_Mux_8_i31_4_lut (.A(n52593), .B(\next_i2c_device_driver_state[2] ), 
         .C(\next_i2c_device_driver_state[4] ), .D(n4), .Z(next_data_reg_15__N_362[8])) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam led_data_out_4__I_0_858_Mux_8_i31_4_lut.init = 16'hca0a;
    LUT4 i19763_3_lut_rep_414 (.A(n30434), .B(n30433), .C(n30432), .Z(n52350)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19763_3_lut_rep_414.init = 16'hcaca;
    LUT4 i1_2_lut_rep_274_3_lut_4_lut (.A(resetn), .B(wd_event_active), 
         .C(n53892), .D(resetn_imu_N_1182), .Z(n52210)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(371[14:35])
    defparam i1_2_lut_rep_274_3_lut_4_lut.init = 16'h2000;
    LUT4 i1_2_lut_4_lut_adj_375 (.A(n30434), .B(n30433), .C(n30432), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_4__6__N_624)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_375.init = 16'hca00;
    LUT4 i19759_3_lut_rep_415 (.A(n30430), .B(n30429), .C(n30428), .Z(n52351)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19759_3_lut_rep_415.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_376 (.A(n30430), .B(n30429), .C(n30428), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_4__7__N_618)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_376.init = 16'hca00;
    LUT4 i19751_3_lut_rep_416 (.A(n30422), .B(n30421), .C(n30420), .Z(n52352)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19751_3_lut_rep_416.init = 16'hcaca;
    LUT4 i39524_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52354), 
         .Z(VL53L1X_data_rx_reg_5__2__N_602)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39524_3_lut.init = 16'h5757;
    LUT4 i1_2_lut_4_lut_adj_377 (.A(n30422), .B(n30421), .C(n30420), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_5__1__N_606)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_377.init = 16'hca00;
    LUT4 i39527_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52352), 
         .Z(VL53L1X_data_rx_reg_5__1__N_608)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39527_3_lut.init = 16'h5757;
    CCU2D add_8435_2 (.A0(VL53L1X_osc_cal_val[1]), .B0(VL53L1X_osc_cal_val[0]), 
          .C0(GND_net), .D0(GND_net), .A1(VL53L1X_osc_cal_val[2]), .B1(VL53L1X_osc_cal_val[1]), 
          .C1(GND_net), .D1(GND_net), .COUT(n43967), .S1(next_VL53L1X_measurement_period_31__N_1103[2]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_8435_2.INIT0 = 16'h7000;
    defparam add_8435_2.INIT1 = 16'h5666;
    defparam add_8435_2.INJECT1_0 = "NO";
    defparam add_8435_2.INJECT1_1 = "NO";
    CCU2D add_8268_cout (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n43966), 
          .S0(n17827));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_8268_cout.INIT0 = 16'h0000;
    defparam add_8268_cout.INIT1 = 16'h0000;
    defparam add_8268_cout.INJECT1_0 = "NO";
    defparam add_8268_cout.INJECT1_1 = "NO";
    CCU2D add_8268_16 (.A0(VL53L1X_osc_cal_val[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(VL53L1X_osc_cal_val[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43965), .COUT(n43966), .S0(n17807[17]), 
          .S1(n17807[18]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_8268_16.INIT0 = 16'hfaaa;
    defparam add_8268_16.INIT1 = 16'hfaaa;
    defparam add_8268_16.INJECT1_0 = "NO";
    defparam add_8268_16.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_378 (.A(n34), .B(VL53L1X_measurement_period[7]), .C(VL53L1X_measurement_period[15]), 
         .D(measurement_period_tx_index[0]), .Z(n20_adj_5297)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_378.init = 16'ha088;
    CCU2D add_8268_14 (.A0(VL53L1X_osc_cal_val[14]), .B0(VL53L1X_osc_cal_val[12]), 
          .C0(GND_net), .D0(GND_net), .A1(VL53L1X_osc_cal_val[15]), .B1(VL53L1X_osc_cal_val[13]), 
          .C1(GND_net), .D1(GND_net), .CIN(n43964), .COUT(n43965), .S0(n17807[15]), 
          .S1(n17807[16]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_8268_14.INIT0 = 16'h5666;
    defparam add_8268_14.INIT1 = 16'h5666;
    defparam add_8268_14.INJECT1_0 = "NO";
    defparam add_8268_14.INJECT1_1 = "NO";
    CCU2D add_409_5 (.A0(cal_reg_addr[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(cal_reg_addr[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43784), .COUT(n43785), .S0(next_cal_reg_addr_7__N_1124[3]), 
          .S1(next_cal_reg_addr_7__N_1124[4]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(602[42:66])
    defparam add_409_5.INIT0 = 16'h5aaa;
    defparam add_409_5.INIT1 = 16'h5aaa;
    defparam add_409_5.INJECT1_0 = "NO";
    defparam add_409_5.INJECT1_1 = "NO";
    LUT4 i1_2_lut_adj_379 (.A(data_tx[7]), .B(\next_i2c_device_driver_state[0] ), 
         .Z(n16)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i1_2_lut_adj_379.init = 16'h8888;
    PFUMX i40893 (.BLUT(n52124), .ALUT(n52121), .C0(\next_i2c_device_driver_state[4] ), 
          .Z(next_i2c_state_4__N_386[4]));
    CCU2D add_8268_12 (.A0(VL53L1X_osc_cal_val[12]), .B0(VL53L1X_osc_cal_val[10]), 
          .C0(GND_net), .D0(GND_net), .A1(VL53L1X_osc_cal_val[13]), .B1(VL53L1X_osc_cal_val[11]), 
          .C1(GND_net), .D1(GND_net), .CIN(n43963), .COUT(n43964), .S0(n17807[13]), 
          .S1(n17807[14]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_8268_12.INIT0 = 16'h5666;
    defparam add_8268_12.INIT1 = 16'h5666;
    defparam add_8268_12.INJECT1_0 = "NO";
    defparam add_8268_12.INJECT1_1 = "NO";
    CCU2D add_8268_10 (.A0(VL53L1X_osc_cal_val[10]), .B0(VL53L1X_osc_cal_val[8]), 
          .C0(GND_net), .D0(GND_net), .A1(VL53L1X_osc_cal_val[11]), .B1(VL53L1X_osc_cal_val[9]), 
          .C1(GND_net), .D1(GND_net), .CIN(n43962), .COUT(n43963), .S0(n17807[11]), 
          .S1(n17807[12]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_8268_10.INIT0 = 16'h5666;
    defparam add_8268_10.INIT1 = 16'h5666;
    defparam add_8268_10.INJECT1_0 = "NO";
    defparam add_8268_10.INJECT1_1 = "NO";
    PFUMX i40890 (.BLUT(n52290), .ALUT(n52122), .C0(\next_i2c_device_driver_state[2] ), 
          .Z(n52123));
    CCU2D add_8268_8 (.A0(VL53L1X_osc_cal_val[8]), .B0(VL53L1X_osc_cal_val[6]), 
          .C0(GND_net), .D0(GND_net), .A1(VL53L1X_osc_cal_val[9]), .B1(VL53L1X_osc_cal_val[7]), 
          .C1(GND_net), .D1(GND_net), .CIN(n43961), .COUT(n43962), .S0(n17807[9]), 
          .S1(n17807[10]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_8268_8.INIT0 = 16'h5666;
    defparam add_8268_8.INIT1 = 16'h5666;
    defparam add_8268_8.INJECT1_0 = "NO";
    defparam add_8268_8.INJECT1_1 = "NO";
    CCU2D add_8268_6 (.A0(VL53L1X_osc_cal_val[6]), .B0(VL53L1X_osc_cal_val[4]), 
          .C0(GND_net), .D0(GND_net), .A1(VL53L1X_osc_cal_val[7]), .B1(VL53L1X_osc_cal_val[5]), 
          .C1(GND_net), .D1(GND_net), .CIN(n43960), .COUT(n43961), .S0(n17807[7]), 
          .S1(n17807[8]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_8268_6.INIT0 = 16'h5666;
    defparam add_8268_6.INIT1 = 16'h5666;
    defparam add_8268_6.INJECT1_0 = "NO";
    defparam add_8268_6.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_16 (.A0(count_ms[14]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_ms[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43851), .S0(n44[14]), .S1(n44[15]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(201[41:57])
    defparam sub_10_add_2_16.INIT0 = 16'h5555;
    defparam sub_10_add_2_16.INIT1 = 16'h5555;
    defparam sub_10_add_2_16.INJECT1_0 = "NO";
    defparam sub_10_add_2_16.INJECT1_1 = "NO";
    LUT4 i11363_3_lut (.A(n52380), .B(data_rx[3]), .C(n28247), .Z(VL53L1X_data_rx_reg_7__7__N_472[59])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i11363_3_lut.init = 16'hcaca;
    LUT4 i4_4_lut_rep_535 (.A(n7_adj_5271), .B(n7250), .C(\next_i2c_device_driver_state[0] ), 
         .D(n52210), .Z(sys_clk_enable_123)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i4_4_lut_rep_535.init = 16'h8000;
    LUT4 i39530_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(\VL53L1X_data_rx_reg[5] [0]), 
         .Z(VL53L1X_data_rx_reg_5__0__N_614)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39530_3_lut.init = 16'h5757;
    LUT4 i23383_3_lut (.A(cal_reg_addr[1]), .B(data_reg[1]), .C(\next_i2c_device_driver_state[0] ), 
         .Z(n34032)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i23383_3_lut.init = 16'hcaca;
    LUT4 i39533_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52351), 
         .Z(VL53L1X_data_rx_reg_4__7__N_620)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39533_3_lut.init = 16'h5757;
    CCU2D add_8268_4 (.A0(VL53L1X_osc_cal_val[4]), .B0(VL53L1X_osc_cal_val[2]), 
          .C0(GND_net), .D0(GND_net), .A1(VL53L1X_osc_cal_val[5]), .B1(VL53L1X_osc_cal_val[3]), 
          .C1(GND_net), .D1(GND_net), .CIN(n43959), .COUT(n43960), .S0(n17807[5]), 
          .S1(n17807[6]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_8268_4.INIT0 = 16'h5666;
    defparam add_8268_4.INIT1 = 16'h5666;
    defparam add_8268_4.INJECT1_0 = "NO";
    defparam add_8268_4.INJECT1_1 = "NO";
    LUT4 i11332_3_lut (.A(n52381), .B(data_rx[4]), .C(n28247), .Z(VL53L1X_data_rx_reg_7__7__N_472[60])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i11332_3_lut.init = 16'hcaca;
    LUT4 i11315_3_lut (.A(n52384), .B(data_rx[5]), .C(n28247), .Z(VL53L1X_data_rx_reg_7__7__N_472[61])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i11315_3_lut.init = 16'hcaca;
    LUT4 i37_else_4_lut (.A(n53892), .B(\next_i2c_device_driver_state[0] ), 
         .C(\next_i2c_device_driver_state[3] ), .D(\next_i2c_device_driver_state[4] ), 
         .Z(n52513)) /* synthesis lut_function=(A (B (D)+!B !(C))+!A !(C (D))) */ ;
    defparam i37_else_4_lut.init = 16'h8f57;
    CCU2D add_8268_2 (.A0(VL53L1X_osc_cal_val[2]), .B0(VL53L1X_osc_cal_val[0]), 
          .C0(GND_net), .D0(GND_net), .A1(VL53L1X_osc_cal_val[3]), .B1(VL53L1X_osc_cal_val[1]), 
          .C1(GND_net), .D1(GND_net), .COUT(n43959), .S1(n17807[4]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_8268_2.INIT0 = 16'h7000;
    defparam add_8268_2.INIT1 = 16'h5666;
    defparam add_8268_2.INJECT1_0 = "NO";
    defparam add_8268_2.INJECT1_1 = "NO";
    PFUMX i40865 (.BLUT(n52086), .ALUT(n49433), .C0(\next_i2c_device_driver_state[3] ), 
          .Z(n52087));
    LUT4 i20005_1_lut (.A(count_ms[15]), .Z(n30677)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam i20005_1_lut.init = 16'h5555;
    LUT4 i11232_2_lut (.A(count_sys_clk_for_ms[16]), .B(n7654[7]), .Z(n21625)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam i11232_2_lut.init = 16'h8888;
    LUT4 i39536_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52350), 
         .Z(VL53L1X_data_rx_reg_4__6__N_626)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39536_3_lut.init = 16'h5757;
    L6MUX21 led_data_out_4__I_0_860_Mux_0_i31 (.D0(n49510), .D1(n49512), 
            .SD(n49571), .Z(next_i2c_state_4__N_386[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;
    PFUMX i38717 (.BLUT(n49511), .ALUT(n30_adj_5320), .C0(\next_i2c_device_driver_state[4] ), 
          .Z(n49512));
    PFUMX i40858 (.BLUT(n52077), .ALUT(n52076), .C0(measurement_period_tx_index[0]), 
          .Z(n52078));
    LUT4 i39539_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52348), 
         .Z(VL53L1X_data_rx_reg_4__5__N_632)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39539_3_lut.init = 16'h5757;
    LUT4 i39542_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52347), 
         .Z(VL53L1X_data_rx_reg_4__4__N_638)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39542_3_lut.init = 16'h5757;
    CCU2D add_8527_18 (.A0(n25[21]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n25[22]), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n43956), 
          .S0(next_VL53L1X_measurement_period_31__N_1103[21]), .S1(next_VL53L1X_measurement_period_31__N_1103[22]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_8527_18.INIT0 = 16'h5aaa;
    defparam add_8527_18.INIT1 = 16'h5aaa;
    defparam add_8527_18.INJECT1_0 = "NO";
    defparam add_8527_18.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_14 (.A0(count_ms[12]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_ms[13]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43850), .COUT(n43851), .S0(n44[12]), .S1(n44[13]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(201[41:57])
    defparam sub_10_add_2_14.INIT0 = 16'h5555;
    defparam sub_10_add_2_14.INIT1 = 16'h5555;
    defparam sub_10_add_2_14.INJECT1_0 = "NO";
    defparam sub_10_add_2_14.INJECT1_1 = "NO";
    PFUMX led_data_out_4__I_0_859_Mux_6_i31 (.BLUT(n14), .ALUT(n15_adj_5291), 
          .C0(n49665), .Z(next_data_tx_7__N_378[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;
    LUT4 i39545_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52346), 
         .Z(VL53L1X_data_rx_reg_4__3__N_644)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39545_3_lut.init = 16'h5757;
    LUT4 i19747_3_lut_rep_418 (.A(n30418), .B(n30417), .C(n30416), .Z(n52354)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19747_3_lut_rep_418.init = 16'hcaca;
    PFUMX i40835 (.BLUT(n52041), .ALUT(n52040), .C0(\next_i2c_device_driver_state[4] ), 
          .Z(n52042));
    LUT4 i1_2_lut_4_lut_adj_380 (.A(n30418), .B(n30417), .C(n30416), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_5__2__N_600)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_380.init = 16'hca00;
    PFUMX led_data_out_4__I_0_859_Mux_4_i31 (.BLUT(n23405), .ALUT(n23389), 
          .C0(\next_i2c_device_driver_state[4] ), .Z(next_data_tx_7__N_378[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;
    CCU2D add_8527_16 (.A0(n25[19]), .B0(VL53L1X_osc_cal_val[14]), .C0(GND_net), 
          .D0(GND_net), .A1(n25[20]), .B1(VL53L1X_osc_cal_val[15]), .C1(GND_net), 
          .D1(GND_net), .CIN(n43955), .COUT(n43956), .S0(next_VL53L1X_measurement_period_31__N_1103[19]), 
          .S1(next_VL53L1X_measurement_period_31__N_1103[20]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_8527_16.INIT0 = 16'h5666;
    defparam add_8527_16.INIT1 = 16'h5666;
    defparam add_8527_16.INJECT1_0 = "NO";
    defparam add_8527_16.INJECT1_1 = "NO";
    LUT4 i26961_4_lut (.A(cal_reg_addr[6]), .B(n37517), .C(data_reg[6]), 
         .D(\next_i2c_device_driver_state[0] ), .Z(n14_adj_5296)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam i26961_4_lut.init = 16'hc088;
    LUT4 i39548_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52345), 
         .Z(VL53L1X_data_rx_reg_4__2__N_650)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39548_3_lut.init = 16'h5757;
    CCU2D add_8527_14 (.A0(n25[17]), .B0(VL53L1X_osc_cal_val[12]), .C0(GND_net), 
          .D0(GND_net), .A1(n25[18]), .B1(VL53L1X_osc_cal_val[13]), .C1(GND_net), 
          .D1(GND_net), .CIN(n43954), .COUT(n43955), .S0(next_VL53L1X_measurement_period_31__N_1103[17]), 
          .S1(next_VL53L1X_measurement_period_31__N_1103[18]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_8527_14.INIT0 = 16'h5666;
    defparam add_8527_14.INIT1 = 16'h5666;
    defparam add_8527_14.INJECT1_0 = "NO";
    defparam add_8527_14.INJECT1_1 = "NO";
    LUT4 i26853_4_lut (.A(cal_reg_addr[3]), .B(n37517), .C(data_reg[3]), 
         .D(\next_i2c_device_driver_state[0] ), .Z(n14_adj_5295)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam i26853_4_lut.init = 16'hc088;
    LUT4 i39551_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52344), 
         .Z(VL53L1X_data_rx_reg_4__1__N_656)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39551_3_lut.init = 16'h5757;
    LUT4 i39554_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52343), 
         .Z(VL53L1X_data_rx_reg_4__0__N_662)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39554_3_lut.init = 16'h5757;
    CCU2D add_8527_12 (.A0(n25[15]), .B0(VL53L1X_osc_cal_val[10]), .C0(GND_net), 
          .D0(GND_net), .A1(n25[16]), .B1(VL53L1X_osc_cal_val[11]), .C1(GND_net), 
          .D1(GND_net), .CIN(n43953), .COUT(n43954), .S0(next_VL53L1X_measurement_period_31__N_1103[15]), 
          .S1(next_VL53L1X_measurement_period_31__N_1103[16]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_8527_12.INIT0 = 16'h5666;
    defparam add_8527_12.INIT1 = 16'h5666;
    defparam add_8527_12.INJECT1_0 = "NO";
    defparam add_8527_12.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_12 (.A0(count_ms[10]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_ms[11]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43849), .COUT(n43850), .S0(n44[10]), .S1(n44[11]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(201[41:57])
    defparam sub_10_add_2_12.INIT0 = 16'h5555;
    defparam sub_10_add_2_12.INIT1 = 16'h5555;
    defparam sub_10_add_2_12.INJECT1_0 = "NO";
    defparam sub_10_add_2_12.INJECT1_1 = "NO";
    LUT4 n33838_bdd_4_lut_40182_4_lut (.A(n52283), .B(\next_i2c_device_driver_return_state[0] ), 
         .C(\next_i2c_device_driver_state[4] ), .D(\next_i2c_device_driver_state[0] ), 
         .Z(n50826)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B+!((D)+!C))) */ ;
    defparam n33838_bdd_4_lut_40182_4_lut.init = 16'hc4f4;
    LUT4 i19743_3_lut_rep_421 (.A(n30414), .B(n30413), .C(n30412), .Z(n52357)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19743_3_lut_rep_421.init = 16'hcaca;
    LUT4 data_tx_1__bdd_4_lut_4_lut (.A(n52283), .B(\next_i2c_device_driver_state[3] ), 
         .C(n14_adj_5335), .D(data_tx[1]), .Z(n52135)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;
    defparam data_tx_1__bdd_4_lut_4_lut.init = 16'hd1c0;
    LUT4 i1_2_lut_4_lut_adj_381 (.A(n30414), .B(n30413), .C(n30412), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_5__3__N_594)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_381.init = 16'hca00;
    LUT4 n33838_bdd_4_lut_4_lut (.A(n52283), .B(\next_i2c_device_driver_state[3] ), 
         .C(n51024), .D(data_tx[0]), .Z(n52157)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;
    defparam n33838_bdd_4_lut_4_lut.init = 16'hd1c0;
    LUT4 i19739_3_lut_rep_422 (.A(n30410), .B(n30409), .C(n30408), .Z(n52358)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19739_3_lut_rep_422.init = 16'hcaca;
    LUT4 i38682_4_lut_4_lut (.A(n52283), .B(\next_i2c_device_driver_return_state[1] ), 
         .C(\next_i2c_device_driver_state[3] ), .D(n14_adj_5270), .Z(n49477)) /* synthesis lut_function=(A (C (D))+!A (B ((D)+!C)+!B (C (D)))) */ ;
    defparam i38682_4_lut_4_lut.init = 16'hf404;
    CCU2D add_8527_10 (.A0(n25[13]), .B0(VL53L1X_osc_cal_val[8]), .C0(GND_net), 
          .D0(GND_net), .A1(n25[14]), .B1(VL53L1X_osc_cal_val[9]), .C1(GND_net), 
          .D1(GND_net), .CIN(n43952), .COUT(n43953), .S0(next_VL53L1X_measurement_period_31__N_1103[13]), 
          .S1(next_VL53L1X_measurement_period_31__N_1103[14]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_8527_10.INIT0 = 16'h5666;
    defparam add_8527_10.INIT1 = 16'h5666;
    defparam add_8527_10.INJECT1_0 = "NO";
    defparam add_8527_10.INJECT1_1 = "NO";
    LUT4 i1_2_lut_4_lut_adj_382 (.A(n30410), .B(n30409), .C(n30408), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_5__4__N_588)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_382.init = 16'hca00;
    LUT4 i11282_3_lut (.A(n52386), .B(data_rx[6]), .C(n28247), .Z(VL53L1X_data_rx_reg_7__7__N_472[62])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i11282_3_lut.init = 16'hcaca;
    LUT4 i39557_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52340), 
         .Z(VL53L1X_data_rx_reg_1__7__N_684)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39557_3_lut.init = 16'h5757;
    LUT4 i39907_4_lut (.A(n7250), .B(n27), .C(n52296), .D(n7246), .Z(sys_clk_enable_254)) /* synthesis lut_function=(!(A+(B (C+!(D))+!B (C (D))))) */ ;
    defparam i39907_4_lut.init = 16'h0511;
    LUT4 i11260_3_lut (.A(\VL53L1X_data_rx_reg[7] [7]), .B(data_rx[7]), 
         .C(n28247), .Z(VL53L1X_data_rx_reg_7__7__N_472[63])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i11260_3_lut.init = 16'hcaca;
    CCU2D add_8527_8 (.A0(n25[11]), .B0(VL53L1X_osc_cal_val[6]), .C0(GND_net), 
          .D0(GND_net), .A1(n25[12]), .B1(VL53L1X_osc_cal_val[7]), .C1(GND_net), 
          .D1(GND_net), .CIN(n43951), .COUT(n43952), .S0(next_VL53L1X_measurement_period_31__N_1103[11]), 
          .S1(next_VL53L1X_measurement_period_31__N_1103[12]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_8527_8.INIT0 = 16'h5666;
    defparam add_8527_8.INIT1 = 16'h5666;
    defparam add_8527_8.INJECT1_0 = "NO";
    defparam add_8527_8.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_10 (.A0(count_ms[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_ms[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43848), .COUT(n43849), .S0(count_ms_15__N_894[8]), 
          .S1(count_ms_15__N_894[9]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(201[41:57])
    defparam sub_10_add_2_10.INIT0 = 16'h5555;
    defparam sub_10_add_2_10.INIT1 = 16'h5555;
    defparam sub_10_add_2_10.INJECT1_0 = "NO";
    defparam sub_10_add_2_10.INJECT1_1 = "NO";
    LUT4 i32_3_lut (.A(\next_i2c_device_driver_state[0] ), .B(n7234), .C(n7240), 
         .Z(n27)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;
    defparam i32_3_lut.init = 16'h3a3a;
    LUT4 mux_5289_i2_4_lut (.A(n52203), .B(n6), .C(n7246), .D(n52296), 
         .Z(n13181[1])) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (B+((D)+!C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam mux_5289_i2_4_lut.init = 16'h0a3a;
    LUT4 i39578_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52333), 
         .Z(VL53L1X_data_rx_reg_1__0__N_726)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39578_3_lut.init = 16'h5757;
    CCU2D add_8527_6 (.A0(n25[9]), .B0(VL53L1X_osc_cal_val[4]), .C0(GND_net), 
          .D0(GND_net), .A1(n25[10]), .B1(VL53L1X_osc_cal_val[5]), .C1(GND_net), 
          .D1(GND_net), .CIN(n43950), .COUT(n43951), .S0(next_VL53L1X_measurement_period_31__N_1103[9]), 
          .S1(next_VL53L1X_measurement_period_31__N_1103[10]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_8527_6.INIT0 = 16'h5666;
    defparam add_8527_6.INIT1 = 16'h5666;
    defparam add_8527_6.INJECT1_0 = "NO";
    defparam add_8527_6.INJECT1_1 = "NO";
    LUT4 i25648_4_lut (.A(n52314), .B(n53890), .C(n30), .D(\next_i2c_device_driver_state[4] ), 
         .Z(next_target_read_count[0])) /* synthesis lut_function=(A (B+!(C (D)))+!A (B+!(C+!(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(395[14] 871[12])
    defparam i25648_4_lut.init = 16'hcfee;
    LUT4 i39445_4_lut (.A(n52303), .B(n53892), .C(n52246), .D(n7250), 
         .Z(n49101)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam i39445_4_lut.init = 16'h2000;
    CCU2D add_8527_4 (.A0(n25[7]), .B0(VL53L1X_osc_cal_val[2]), .C0(GND_net), 
          .D0(GND_net), .A1(n25[8]), .B1(VL53L1X_osc_cal_val[3]), .C1(GND_net), 
          .D1(GND_net), .CIN(n43949), .COUT(n43950), .S0(next_VL53L1X_measurement_period_31__N_1103[7]), 
          .S1(next_VL53L1X_measurement_period_31__N_1103[8]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_8527_4.INIT0 = 16'h5666;
    defparam add_8527_4.INIT1 = 16'h5666;
    defparam add_8527_4.INJECT1_0 = "NO";
    defparam add_8527_4.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_8 (.A0(count_ms[6]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_ms[7]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43847), .COUT(n43848), .S0(count_ms_15__N_894[6]), 
          .S1(count_ms_15__N_894[7]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(201[41:57])
    defparam sub_10_add_2_8.INIT0 = 16'h5555;
    defparam sub_10_add_2_8.INIT1 = 16'h5555;
    defparam sub_10_add_2_8.INJECT1_0 = "NO";
    defparam sub_10_add_2_8.INJECT1_1 = "NO";
    LUT4 mux_3485_i1_4_lut (.A(n53), .B(\next_i2c_device_driver_state[3] ), 
         .C(n6972), .D(n52447), .Z(n6915[0])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(395[14] 871[12])
    defparam mux_3485_i1_4_lut.init = 16'hc5c0;
    LUT4 i12_3_lut (.A(valid_strobe_enable), .B(throttle_controller_active), 
         .C(next_imu_data_valid), .Z(valid_strobe_N_1132)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(299[14] 304[12])
    defparam i12_3_lut.init = 16'h3a3a;
    LUT4 VL53L1X_data_rx_reg_index_i1_i2_3_lut (.A(n52446), .B(n52447), 
         .C(one_byte_ready), .Z(n23[1])) /* synthesis lut_function=(!(A (B (C))+!A !(B (C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(229[14] 230[75])
    defparam VL53L1X_data_rx_reg_index_i1_i2_3_lut.init = 16'h6a6a;
    CCU2D add_8527_2 (.A0(n25[5]), .B0(VL53L1X_osc_cal_val[0]), .C0(GND_net), 
          .D0(GND_net), .A1(n25[6]), .B1(VL53L1X_osc_cal_val[1]), .C1(GND_net), 
          .D1(GND_net), .COUT(n43949), .S1(next_VL53L1X_measurement_period_31__N_1103[6]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(705[57:84])
    defparam add_8527_2.INIT0 = 16'h7000;
    defparam add_8527_2.INIT1 = 16'h5666;
    defparam add_8527_2.INJECT1_0 = "NO";
    defparam add_8527_2.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_6 (.A0(count_ms[4]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_ms[5]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43846), .COUT(n43847), .S0(count_ms_15__N_894[4]), 
          .S1(count_ms_15__N_894[5]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(201[41:57])
    defparam sub_10_add_2_6.INIT0 = 16'h5555;
    defparam sub_10_add_2_6.INIT1 = 16'h5555;
    defparam sub_10_add_2_6.INJECT1_0 = "NO";
    defparam sub_10_add_2_6.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_4 (.A0(count_ms[2]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_ms[3]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43845), .COUT(n43846), .S0(count_ms_15__N_894[2]), 
          .S1(n44[3]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(201[41:57])
    defparam sub_10_add_2_4.INIT0 = 16'h5555;
    defparam sub_10_add_2_4.INIT1 = 16'h5555;
    defparam sub_10_add_2_4.INJECT1_0 = "NO";
    defparam sub_10_add_2_4.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_2 (.A0(count_ms[0]), .B0(count_ms[15]), .C0(GND_net), 
          .D0(GND_net), .A1(count_ms[1]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n43845), .S1(count_ms_15__N_894[1]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(201[41:57])
    defparam sub_10_add_2_2.INIT0 = 16'h1000;
    defparam sub_10_add_2_2.INIT1 = 16'h5555;
    defparam sub_10_add_2_2.INJECT1_0 = "NO";
    defparam sub_10_add_2_2.INJECT1_1 = "NO";
    CCU2D add_409_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(cal_reg_addr[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n43783), .S1(next_cal_reg_addr_7__N_1124[0]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(602[42:66])
    defparam add_409_1.INIT0 = 16'hF000;
    defparam add_409_1.INIT1 = 16'h5555;
    defparam add_409_1.INJECT1_0 = "NO";
    defparam add_409_1.INJECT1_1 = "NO";
    LUT4 i1_4_lut_4_lut_then_3_lut_adj_383 (.A(\next_i2c_device_driver_state[3] ), 
         .B(\next_i2c_device_driver_state[0] ), .C(next_i2c_state_4__N_1050[0]), 
         .Z(n52508)) /* synthesis lut_function=((B+!(C))+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i1_4_lut_4_lut_then_3_lut_adj_383.init = 16'hdfdf;
    L6MUX21 i38714 (.D0(n49507), .D1(n49508), .SD(\next_i2c_device_driver_state[4] ), 
            .Z(next_i2c_state_4__N_386[1]));
    LUT4 i39560_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52339), 
         .Z(VL53L1X_data_rx_reg_1__6__N_690)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39560_3_lut.init = 16'h5757;
    LUT4 i26488_2_lut (.A(data_tx[0]), .B(\next_i2c_device_driver_state[0] ), 
         .Z(n19_adj_5319)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam i26488_2_lut.init = 16'h8888;
    LUT4 i39950_2_lut_rep_536 (.A(resetn), .B(wd_event_active), .C(n52306), 
         .D(\i2c_top_debug[1] ), .Z(n53890)) /* synthesis lut_function=((B+!(C+(D)))+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(371[14:35])
    defparam i39950_2_lut_rep_536.init = 16'hdddf;
    LUT4 i39563_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52338), 
         .Z(VL53L1X_data_rx_reg_1__5__N_696)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39563_3_lut.init = 16'h5757;
    LUT4 i39581_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52332), 
         .Z(VL53L1X_data_rx_reg_0__7__N_732)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39581_3_lut.init = 16'h5757;
    PFUMX i40172 (.BLUT(n51006), .ALUT(n51005), .C0(\next_i2c_device_driver_state[3] ), 
          .Z(n51007));
    PFUMX i38712 (.BLUT(n7_adj_5325), .ALUT(n22527), .C0(\next_i2c_device_driver_state[3] ), 
          .Z(n49507));
    LUT4 i39584_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52331), 
         .Z(VL53L1X_data_rx_reg_0__6__N_738)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39584_3_lut.init = 16'h5757;
    PFUMX mux_3602_i5 (.BLUT(n13181[4]), .ALUT(n13173[2]), .C0(n7250), 
          .Z(n2485[4]));
    PFUMX mux_3602_i4 (.BLUT(n13181[3]), .ALUT(n13173[1]), .C0(n7250), 
          .Z(n2485[3]));
    CCU2D sub_257_add_2_21 (.A0(master_trigger_count_ms[19]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(master_trigger_count_ms[20]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n43805), .S0(master_trigger_count_ms_20__N_997[19]), 
          .S1(n611[20]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(279[40:72])
    defparam sub_257_add_2_21.INIT0 = 16'h5555;
    defparam sub_257_add_2_21.INIT1 = 16'h5555;
    defparam sub_257_add_2_21.INJECT1_0 = "NO";
    defparam sub_257_add_2_21.INJECT1_1 = "NO";
    LUT4 i39587_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52330), 
         .Z(VL53L1X_data_rx_reg_0__5__N_744)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39587_3_lut.init = 16'h5757;
    LUT4 i39590_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52329), 
         .Z(VL53L1X_data_rx_reg_0__4__N_750)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39590_3_lut.init = 16'h5757;
    CCU2D sub_257_add_2_19 (.A0(master_trigger_count_ms[17]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(master_trigger_count_ms[18]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n43804), .COUT(n43805), 
          .S0(master_trigger_count_ms_20__N_997[17]), .S1(n611[18]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(279[40:72])
    defparam sub_257_add_2_19.INIT0 = 16'h5555;
    defparam sub_257_add_2_19.INIT1 = 16'h5555;
    defparam sub_257_add_2_19.INJECT1_0 = "NO";
    defparam sub_257_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_257_add_2_17 (.A0(master_trigger_count_ms[15]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(master_trigger_count_ms[16]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n43803), .COUT(n43804), 
          .S0(master_trigger_count_ms_20__N_997[15]), .S1(master_trigger_count_ms_20__N_997[16]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(279[40:72])
    defparam sub_257_add_2_17.INIT0 = 16'h5555;
    defparam sub_257_add_2_17.INIT1 = 16'h5555;
    defparam sub_257_add_2_17.INJECT1_0 = "NO";
    defparam sub_257_add_2_17.INJECT1_1 = "NO";
    PFUMX i38713 (.BLUT(n28_adj_5327), .ALUT(n29_adj_5300), .C0(n49625), 
          .Z(n49508));
    LUT4 i19731_3_lut_rep_427 (.A(n30402), .B(n30401), .C(n30400), .Z(n52363)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19731_3_lut_rep_427.init = 16'hcaca;
    LUT4 mux_833_Mux_6_i127_4_lut (.A(n50953), .B(cal_reg_addr[0]), .C(cal_reg_addr[7]), 
         .D(n47344), .Z(n127_adj_5337)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (B+((D)+!C)))) */ ;
    defparam mux_833_Mux_6_i127_4_lut.init = 16'h0a3a;
    LUT4 i1_2_lut_4_lut_adj_384 (.A(n30402), .B(n30401), .C(n30400), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_5__6__N_576)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_384.init = 16'hca00;
    LUT4 i39593_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52324), 
         .Z(VL53L1X_data_rx_reg_0__3__N_756)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39593_3_lut.init = 16'h5757;
    LUT4 i12345_3_lut (.A(n53888), .B(n611[20]), .C(master_trigger_count_ms[20]), 
         .Z(master_trigger_count_ms_20__N_997[20])) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(278[14] 281[12])
    defparam i12345_3_lut.init = 16'hecec;
    LUT4 i6153_1_lut (.A(count_sys_clk_for_ms[16]), .Z(n14054)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam i6153_1_lut.init = 16'h5555;
    LUT4 i19727_3_lut_rep_428 (.A(n30398), .B(n30397), .C(n30396), .Z(n52364)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19727_3_lut_rep_428.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_385 (.A(n30398), .B(n30397), .C(n30396), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_5__7__N_570)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_385.init = 16'hca00;
    PFUMX led_data_out_4__I_0_860_Mux_2_i31 (.BLUT(n14_adj_5288), .ALUT(n15_adj_5280), 
          .C0(n49665), .Z(next_i2c_state_4__N_386[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;
    CCU2D sub_257_add_2_15 (.A0(master_trigger_count_ms[13]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(master_trigger_count_ms[14]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n43802), .COUT(n43803), 
          .S0(n611[13]), .S1(n611[14]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(279[40:72])
    defparam sub_257_add_2_15.INIT0 = 16'h5555;
    defparam sub_257_add_2_15.INIT1 = 16'h5555;
    defparam sub_257_add_2_15.INJECT1_0 = "NO";
    defparam sub_257_add_2_15.INJECT1_1 = "NO";
    LUT4 i17668_4_lut (.A(n52450), .B(\next_i2c_device_driver_return_state[2] ), 
         .C(\next_i2c_device_driver_state[2] ), .D(n28226), .Z(n28220)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C)+!B !((D)+!C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam i17668_4_lut.init = 16'hcafa;
    LUT4 i33208_2_lut (.A(n25[5]), .B(VL53L1X_osc_cal_val[0]), .Z(next_VL53L1X_measurement_period_31__N_1103[5])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i33208_2_lut.init = 16'h6666;
    LUT4 led_data_out_4__I_0_862_Mux_4_i31_4_lut (.A(\next_i2c_device_driver_return_state[4] ), 
         .B(n51007), .C(\next_i2c_device_driver_state[4] ), .D(n25615), 
         .Z(next_return_state_4__N_391[4])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam led_data_out_4__I_0_862_Mux_4_i31_4_lut.init = 16'hc0ca;
    PFUMX i38715 (.BLUT(n1_adj_5338), .ALUT(n3), .C0(n49569), .Z(n49510));
    L6MUX21 i38585 (.D0(n52135), .D1(n53873), .SD(\next_i2c_device_driver_state[4] ), 
            .Z(next_data_tx_7__N_378[1]));
    FD1S3IX i2c_state__i2_rep_538 (.D(next_i2c_state_4__N_386[1]), .CK(sys_clk), 
            .CD(n53891), .Q(n53892)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam i2c_state__i2_rep_538.GSR = "ENABLED";
    PFUMX mux_3602_i8 (.BLUT(n48822), .ALUT(n20052), .C0(n7250), .Z(n2485[7]));
    LUT4 led_data_out_4__I_0_868_Mux_5_i15_4_lut_4_lut (.A(n52271), .B(n52269), 
         .C(\next_i2c_device_driver_state[3] ), .D(next_cal_reg_addr_7__N_1124[5]), 
         .Z(n15_adj_5273)) /* synthesis lut_function=(A (B (C (D)))+!A (B ((D)+!C)+!B !(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam led_data_out_4__I_0_868_Mux_5_i15_4_lut_4_lut.init = 16'hc505;
    LUT4 i19723_3_lut_rep_429 (.A(n30394), .B(n30393), .C(n30392), .Z(n52365)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19723_3_lut_rep_429.init = 16'hcaca;
    LUT4 one_byte_ready_I_0_2_lut_rep_508 (.A(one_byte_ready), .B(rx_from_VL53L1X), 
         .Z(n52444)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[18:51])
    defparam one_byte_ready_I_0_2_lut_rep_508.init = 16'h8888;
    L6MUX21 i61 (.D0(n36), .D1(n27_adj_5339), .SD(i2c_top_debug[2]), .Z(n45689));
    PFUMX i40918 (.BLUT(n52486), .ALUT(n52487), .C0(\next_i2c_device_driver_state[0] ), 
          .Z(n21_adj_5321));
    LUT4 i1_2_lut_rep_282_3_lut_4_lut (.A(one_byte_ready), .B(rx_from_VL53L1X), 
         .C(n52446), .D(VL53L1X_data_rx_reg_index[2]), .Z(n52218)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[18:51])
    defparam i1_2_lut_rep_282_3_lut_4_lut.init = 16'hf7ff;
    LUT4 i1_2_lut_rep_283_3_lut_4_lut (.A(one_byte_ready), .B(rx_from_VL53L1X), 
         .C(n52446), .D(VL53L1X_data_rx_reg_index[2]), .Z(n52219)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[18:51])
    defparam i1_2_lut_rep_283_3_lut_4_lut.init = 16'hfff7;
    LUT4 i1_2_lut_4_lut_adj_386 (.A(n30394), .B(n30393), .C(n30392), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_6__0__N_564)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_386.init = 16'hca00;
    PFUMX i40692 (.BLUT(n51818), .ALUT(n51817), .C0(n7246), .Z(n51819));
    LUT4 i23202_4_lut (.A(n52201), .B(measurement_period_tx_index[0]), .C(\next_i2c_device_driver_state[4] ), 
         .D(n52445), .Z(n33854)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A (B+((D)+!C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i23202_4_lut.init = 16'h0a3a;
    LUT4 i37447_2_lut_rep_320_3_lut (.A(one_byte_ready), .B(rx_from_VL53L1X), 
         .C(VL53L1X_data_rx_reg_index[2]), .Z(n52256)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[18:51])
    defparam i37447_2_lut_rep_320_3_lut.init = 16'h8080;
    CCU2D sub_257_add_2_13 (.A0(master_trigger_count_ms[11]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(master_trigger_count_ms[12]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n43801), .COUT(n43802), 
          .S0(master_trigger_count_ms_20__N_997[11]), .S1(master_trigger_count_ms_20__N_997[12]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(279[40:72])
    defparam sub_257_add_2_13.INIT0 = 16'h5555;
    defparam sub_257_add_2_13.INIT1 = 16'h5555;
    defparam sub_257_add_2_13.INJECT1_0 = "NO";
    defparam sub_257_add_2_13.INJECT1_1 = "NO";
    LUT4 i18924_2_lut_rep_267 (.A(n7234), .B(n7240), .Z(n52203)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam i18924_2_lut_rep_267.init = 16'h8888;
    PFUMX i7 (.BLUT(n14_adj_5340), .ALUT(n6_adj_5313), .C0(n49665), .Z(next_data_reg_15__N_362[4]));
    LUT4 i19719_3_lut_rep_430 (.A(n30390), .B(n30389), .C(n30388), .Z(n52366)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19719_3_lut_rep_430.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_387 (.A(n30390), .B(n30389), .C(n30388), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_6__1__N_558)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_387.init = 16'hca00;
    LUT4 i1_2_lut_rep_509 (.A(measurement_period_tx_index[1]), .B(measurement_period_tx_index[2]), 
         .Z(n52445)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam i1_2_lut_rep_509.init = 16'heeee;
    PFUMX i40139 (.BLUT(n50952), .ALUT(n50951), .C0(cal_reg_addr[6]), 
          .Z(n50953));
    PFUMX i48 (.BLUT(n53877), .ALUT(n28_adj_5285), .C0(\next_i2c_device_driver_state[4] ), 
          .Z(next_data_tx_7__N_378[7]));
    LUT4 i39783_2_lut_3_lut (.A(measurement_period_tx_index[1]), .B(measurement_period_tx_index[2]), 
         .C(\next_i2c_device_driver_state[0] ), .Z(n34)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam i39783_2_lut_3_lut.init = 16'h0101;
    CCU2D sub_257_add_2_11 (.A0(master_trigger_count_ms[9]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(master_trigger_count_ms[10]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n43800), .COUT(n43801), 
          .S0(n611[9]), .S1(n611[10]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(279[40:72])
    defparam sub_257_add_2_11.INIT0 = 16'h5555;
    defparam sub_257_add_2_11.INIT1 = 16'h5555;
    defparam sub_257_add_2_11.INJECT1_0 = "NO";
    defparam sub_257_add_2_11.INJECT1_1 = "NO";
    PFUMX i48_adj_388 (.BLUT(n53879), .ALUT(n28_adj_5282), .C0(\next_i2c_device_driver_state[4] ), 
          .Z(next_data_tx_7__N_378[3]));
    FD1S3IX data_tx__i1 (.D(next_data_tx_7__N_378[1]), .CK(sys_clk), .CD(n52212), 
            .Q(data_tx[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam data_tx__i1.GSR = "ENABLED";
    LUT4 i27164_2_lut_3_lut (.A(\next_i2c_device_driver_state[0] ), .B(\next_i2c_device_driver_return_state[1] ), 
         .C(n53892), .Z(n13)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam i27164_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i19715_3_lut_rep_431 (.A(n30386), .B(n30385), .C(n30384), .Z(n52367)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19715_3_lut_rep_431.init = 16'hcaca;
    LUT4 led_data_out_4__I_0_862_Mux_1_i21_3_lut_3_lut_3_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(\next_i2c_device_driver_return_state[1] ), .C(n53892), .Z(n21_adj_5302)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam led_data_out_4__I_0_862_Mux_1_i21_3_lut_3_lut_3_lut.init = 16'h5858;
    LUT4 i1_2_lut_4_lut_adj_389 (.A(n30386), .B(n30385), .C(n30384), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_6__2__N_552)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_389.init = 16'hca00;
    CCU2D sub_257_add_2_9 (.A0(master_trigger_count_ms[7]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(master_trigger_count_ms[8]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n43799), .COUT(n43800), 
          .S0(master_trigger_count_ms_20__N_997[7]), .S1(n611[8]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(279[40:72])
    defparam sub_257_add_2_9.INIT0 = 16'h5555;
    defparam sub_257_add_2_9.INIT1 = 16'h5555;
    defparam sub_257_add_2_9.INJECT1_0 = "NO";
    defparam sub_257_add_2_9.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_adj_390 (.A(\next_i2c_device_driver_state[0] ), .B(\next_i2c_device_driver_return_state[1] ), 
         .C(next_i2c_state_4__N_1050[0]), .Z(n11_adj_5331)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam i1_2_lut_3_lut_adj_390.init = 16'h8080;
    LUT4 led_data_out_4__I_0_868_Mux_3_i15_4_lut_4_lut (.A(n52271), .B(n52269), 
         .C(\next_i2c_device_driver_state[3] ), .D(next_cal_reg_addr_7__N_1124[3]), 
         .Z(n15_adj_5274)) /* synthesis lut_function=(A (B (C (D)))+!A (B ((D)+!C)+!B !(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam led_data_out_4__I_0_868_Mux_3_i15_4_lut_4_lut.init = 16'hc505;
    LUT4 i19948_3_lut_rep_510 (.A(n30619), .B(n30618), .C(n30617), .Z(n52446)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(229[14] 230[75])
    defparam i19948_3_lut_rep_510.init = 16'hcaca;
    LUT4 led_data_out_4__I_0_868_Mux_2_i15_4_lut_4_lut (.A(n52271), .B(n52269), 
         .C(\next_i2c_device_driver_state[3] ), .D(next_cal_reg_addr_7__N_1124[2]), 
         .Z(n15_adj_5275)) /* synthesis lut_function=(A (B (C (D)))+!A (B ((D)+!C)+!B !(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam led_data_out_4__I_0_868_Mux_2_i15_4_lut_4_lut.init = 16'hc505;
    LUT4 i19711_3_lut_rep_432 (.A(n30382), .B(n30381), .C(n30380), .Z(n52368)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19711_3_lut_rep_432.init = 16'hcaca;
    LUT4 i1_2_lut_rep_356_4_lut (.A(n30619), .B(n30618), .C(n30617), .D(n52447), 
         .Z(n52292)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (((D)+!C)+!B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(229[14] 230[75])
    defparam i1_2_lut_rep_356_4_lut.init = 16'hff35;
    LUT4 i19659_3_lut_rep_511 (.A(n30330), .B(n30329), .C(n30328), .Z(n52447)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(229[14] 230[75])
    defparam i19659_3_lut_rep_511.init = 16'hcaca;
    LUT4 i8566_2_lut_4_lut (.A(n30330), .B(n30329), .C(n30328), .D(one_byte_ready), 
         .Z(n23[0])) /* synthesis lut_function=(!(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B !(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(229[14] 230[75])
    defparam i8566_2_lut_4_lut.init = 16'h35ca;
    LUT4 i39443_2_lut_rep_512 (.A(resetn_VL53L1X_buffer), .B(resetn), .Z(n52448)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i39443_2_lut_rep_512.init = 16'h7777;
    LUT4 i1_2_lut_4_lut_adj_391 (.A(n30382), .B(n30381), .C(n30380), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_6__3__N_546)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_391.init = 16'hca00;
    LUT4 i39455_3_lut_4_lut (.A(resetn_VL53L1X_buffer), .B(resetn), .C(next_VL53L1X_data_rx_reg_index[1]), 
         .D(n48780), .Z(VL53L1X_data_rx_reg_index_5__N_460)) /* synthesis lut_function=(!(A (B (C+(D))))) */ ;
    defparam i39455_3_lut_4_lut.init = 16'h777f;
    LUT4 i19707_3_lut_rep_433 (.A(n30378), .B(n30377), .C(n30376), .Z(n52369)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19707_3_lut_rep_433.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_392 (.A(n30378), .B(n30377), .C(n30376), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_6__4__N_540)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_392.init = 16'hca00;
    LUT4 i39453_3_lut_4_lut (.A(resetn_VL53L1X_buffer), .B(resetn), .C(next_VL53L1X_data_rx_reg_index[2]), 
         .D(n48780), .Z(VL53L1X_data_rx_reg_index_5__N_457)) /* synthesis lut_function=(!(A (B (C+(D))))) */ ;
    defparam i39453_3_lut_4_lut.init = 16'h777f;
    LUT4 i19703_3_lut_rep_434 (.A(n30374), .B(n30373), .C(n30372), .Z(n52370)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19703_3_lut_rep_434.init = 16'hcaca;
    LUT4 VL53L1X_data_rx_reg_index_5__N_427_I_0_749_3_lut_3_lut_4_lut (.A(resetn_VL53L1X_buffer), 
         .B(resetn), .C(next_VL53L1X_data_rx_reg_index[1]), .D(n48780), 
         .Z(VL53L1X_data_rx_reg_index_5__N_442)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam VL53L1X_data_rx_reg_index_5__N_427_I_0_749_3_lut_3_lut_4_lut.init = 16'h0080;
    LUT4 VL53L1X_data_rx_reg_index_5__N_427_I_0_748_3_lut_3_lut_4_lut (.A(resetn_VL53L1X_buffer), 
         .B(resetn), .C(next_VL53L1X_data_rx_reg_index[2]), .D(n48780), 
         .Z(VL53L1X_data_rx_reg_index_5__N_439)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam VL53L1X_data_rx_reg_index_5__N_427_I_0_748_3_lut_3_lut_4_lut.init = 16'h0080;
    LUT4 n6_bdd_2_lut_3_lut (.A(n7234), .B(n7240), .C(is_2_byte_reg), 
         .Z(n51818)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam n6_bdd_2_lut_3_lut.init = 16'hf8f8;
    LUT4 i27338_2_lut_rep_513 (.A(\next_i2c_device_driver_state[0] ), .B(n53892), 
         .Z(n52449)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i27338_2_lut_rep_513.init = 16'heeee;
    LUT4 i1_2_lut_4_lut_adj_393 (.A(n30374), .B(n30373), .C(n30372), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_6__5__N_534)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_393.init = 16'hca00;
    LUT4 i5_1_lut_rep_354_2_lut (.A(\next_i2c_device_driver_state[0] ), .B(n53892), 
         .Z(n52290)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i5_1_lut_rep_354_2_lut.init = 16'h1111;
    LUT4 i39596_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52322), 
         .Z(VL53L1X_data_rx_reg_0__2__N_762)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39596_3_lut.init = 16'h5757;
    LUT4 i1_3_lut_3_lut_4_lut_adj_394 (.A(\next_i2c_device_driver_state[0] ), 
         .B(n53892), .C(\next_i2c_device_driver_return_state[3] ), .D(\next_i2c_device_driver_state[2] ), 
         .Z(n29)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_3_lut_3_lut_4_lut_adj_394.init = 16'hf0ee;
    LUT4 next_i2c_device_driver_state_4__bdd_3_lut_40087_3_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n53892), .C(target_read_count[1]), .D(\next_i2c_device_driver_state[2] ), 
         .Z(n50877)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+(D)))) */ ;
    defparam next_i2c_device_driver_state_4__bdd_3_lut_40087_3_lut_4_lut.init = 16'hf1f0;
    PFUMX led_data_out_4__I_0_859_Mux_2_i31 (.BLUT(n53876), .ALUT(n22284), 
          .C0(\next_i2c_device_driver_state[4] ), .Z(next_data_tx_7__N_378[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;
    LUT4 i23_3_lut_3_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), .B(n53892), 
         .C(\next_i2c_device_driver_state[2] ), .D(\next_i2c_device_driver_state[3] ), 
         .Z(n17_adj_5342)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B (C (D)+!C !(D)))) */ ;
    defparam i23_3_lut_3_lut_4_lut.init = 16'hf0ef;
    LUT4 i39914_2_lut_rep_334_3_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n53892), .C(next_VL53L1X_firm_rdy[0]), .Z(n52270)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam i39914_2_lut_rep_334_3_lut.init = 16'h0101;
    LUT4 i1_2_lut_rep_335_2_lut_3_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n53892), .C(\next_i2c_device_driver_state[2] ), .Z(n52271)) /* synthesis lut_function=(A+(B+!(C))) */ ;
    defparam i1_2_lut_rep_335_2_lut_3_lut.init = 16'hefef;
    PFUMX mux_833_Mux_6_i255 (.BLUT(n125), .ALUT(n127_adj_5337), .C0(n49535), 
          .Z(next_data_tx_7__N_1032_c[6]));
    LUT4 n6_bdd_3_lut_40171_4_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n53892), .C(\next_i2c_device_driver_return_state[4] ), .D(\next_i2c_device_driver_state[2] ), 
         .Z(n51005)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam n6_bdd_3_lut_40171_4_lut.init = 16'hf0ee;
    LUT4 i12_3_lut_3_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), .B(n53892), 
         .C(n48496), .D(\next_i2c_device_driver_state[4] ), .Z(n46519)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam i12_3_lut_3_lut_4_lut.init = 16'hf011;
    LUT4 i39728_2_lut_3_lut (.A(\next_i2c_device_driver_state[0] ), .B(n53892), 
         .C(\next_i2c_device_driver_state[4] ), .Z(n48249)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam i39728_2_lut_3_lut.init = 16'h0101;
    LUT4 i19699_3_lut_rep_435 (.A(n30370), .B(n30369), .C(n30368), .Z(n52371)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19699_3_lut_rep_435.init = 16'hcaca;
    LUT4 i18716_2_lut_rep_514 (.A(\next_i2c_device_driver_state[0] ), .B(n53892), 
         .Z(n52450)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam i18716_2_lut_rep_514.init = 16'h8888;
    LUT4 i1_2_lut_4_lut_adj_395 (.A(n30370), .B(n30369), .C(n30368), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_6__6__N_528)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_395.init = 16'hca00;
    LUT4 i26847_3_lut_3_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n53892), .C(data_reg[3]), .D(\next_i2c_device_driver_state[2] ), 
         .Z(n7_adj_5294)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A ((D)+!C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam i26847_3_lut_3_lut_4_lut.init = 16'h00f8;
    LUT4 i19695_3_lut_rep_436 (.A(n30366), .B(n30365), .C(n30364), .Z(n52372)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19695_3_lut_rep_436.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_396 (.A(n30366), .B(n30365), .C(n30364), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_6__7__N_522)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_396.init = 16'hca00;
    LUT4 i39599_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52321), 
         .Z(VL53L1X_data_rx_reg_0__1__N_768)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39599_3_lut.init = 16'h5757;
    LUT4 i39602_3_lut (.A(resetn), .B(resetn_VL53L1X_buffer), .C(n52320), 
         .Z(VL53L1X_data_rx_reg_0__0__N_774)) /* synthesis lut_function=(!(A (B+(C)))) */ ;
    defparam i39602_3_lut.init = 16'h5757;
    LUT4 i1_2_lut_2_lut_3_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n53892), .C(data_tx[6]), .D(\next_i2c_device_driver_state[2] ), 
         .Z(n7_adj_5290)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam i1_2_lut_2_lut_3_lut_4_lut.init = 16'h0070;
    LUT4 i26920_3_lut_3_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n53892), .C(data_reg[1]), .D(\next_i2c_device_driver_state[2] ), 
         .Z(n7_adj_5293)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A ((D)+!C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam i26920_3_lut_3_lut_4_lut.init = 16'h00f8;
    LUT4 n49433_bdd_3_lut_3_lut_4_lut_3_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n53892), .C(\next_i2c_device_driver_state[2] ), .Z(n52086)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B+!(C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam n49433_bdd_3_lut_3_lut_4_lut_3_lut.init = 16'h1818;
    LUT4 i1_2_lut_rep_347_3_lut (.A(\next_i2c_device_driver_state[0] ), .B(n53892), 
         .C(\next_i2c_device_driver_state[2] ), .Z(n52283)) /* synthesis lut_function=(A (B+(C))+!A (C)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam i1_2_lut_rep_347_3_lut.init = 16'hf8f8;
    LUT4 led_data_out_4__I_0_858_Mux_4_i14_4_lut_4_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n53892), .C(\next_i2c_device_driver_state[2] ), .D(n36072), 
         .Z(n14_adj_5340)) /* synthesis lut_function=(A (B (C)+!B !(C+!(D)))+!A !(B+(C+!(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam led_data_out_4__I_0_858_Mux_4_i14_4_lut_4_lut_4_lut.init = 16'h8380;
    LUT4 next_i2c_device_driver_state_4__bdd_3_lut_40134_3_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n53892), .C(target_read_count[1]), .D(\next_i2c_device_driver_state[2] ), 
         .Z(n50878)) /* synthesis lut_function=(!(A (B (D)+!B ((D)+!C))+!A ((D)+!C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam next_i2c_device_driver_state_4__bdd_3_lut_40134_3_lut_4_lut.init = 16'h00f8;
    PFUMX i40625 (.BLUT(n51725), .ALUT(n51724), .C0(n7250), .Z(n2485[5]));
    LUT4 i1_2_lut_rep_265_2_lut_3_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n53892), .C(\next_i2c_device_driver_return_state[0] ), .D(\next_i2c_device_driver_state[2] ), 
         .Z(n52201)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam i1_2_lut_rep_265_2_lut_3_lut_4_lut.init = 16'h0070;
    PFUMX i40623 (.BLUT(n51722), .ALUT(n51721), .C0(\next_i2c_device_driver_state[2] ), 
          .Z(next_return_state_4__N_391[0]));
    LUT4 n14_bdd_2_lut_3_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n53892), .C(data_reg[4]), .D(\next_i2c_device_driver_state[2] ), 
         .Z(n52041)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam n14_bdd_2_lut_3_lut_4_lut.init = 16'h0070;
    LUT4 i27230_2_lut_2_lut_3_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n53892), .C(data_tx[4]), .Z(n3_adj_5304)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam i27230_2_lut_2_lut_3_lut.init = 16'h7070;
    LUT4 led_data_out_4__I_0_858_Mux_5_i14_4_lut_4_lut_4_lut (.A(\next_i2c_device_driver_state[0] ), 
         .B(n53892), .C(n8_adj_5323), .D(\next_i2c_device_driver_state[2] ), 
         .Z(n14_adj_5277)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A !(B+((D)+!C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam led_data_out_4__I_0_858_Mux_5_i14_4_lut_4_lut_4_lut.init = 16'h8830;
    LUT4 i1_3_lut_4_lut_adj_397 (.A(\next_i2c_device_driver_state[0] ), .B(n53892), 
         .C(n17_adj_5342), .D(\next_i2c_device_driver_state[4] ), .Z(n7250)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam i1_3_lut_4_lut_adj_397.init = 16'hf800;
    CCU2D sub_257_add_2_7 (.A0(master_trigger_count_ms[5]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(master_trigger_count_ms[6]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n43798), .COUT(n43799), 
          .S0(n611[5]), .S1(master_trigger_count_ms_20__N_997[6]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(279[40:72])
    defparam sub_257_add_2_7.INIT0 = 16'h5555;
    defparam sub_257_add_2_7.INIT1 = 16'h5555;
    defparam sub_257_add_2_7.INJECT1_0 = "NO";
    defparam sub_257_add_2_7.INJECT1_1 = "NO";
    PFUMX i40621 (.BLUT(n50826), .ALUT(n51719), .C0(n53892), .Z(n51720));
    PFUMX led_data_out_4__I_0_859_Mux_5_i31 (.BLUT(n53878), .ALUT(n21563), 
          .C0(\next_i2c_device_driver_state[4] ), .Z(next_data_tx_7__N_378[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;
    FD1S3IX data_tx__i2 (.D(next_data_tx_7__N_378[2]), .CK(sys_clk), .CD(n52212), 
            .Q(data_tx[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam data_tx__i2.GSR = "ENABLED";
    FD1S3IX data_tx__i3 (.D(next_data_tx_7__N_378[3]), .CK(sys_clk), .CD(n52212), 
            .Q(data_tx[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam data_tx__i3.GSR = "ENABLED";
    FD1S3IX data_tx__i4 (.D(next_data_tx_7__N_378[4]), .CK(sys_clk), .CD(n52212), 
            .Q(data_tx[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam data_tx__i4.GSR = "ENABLED";
    FD1S3IX data_tx__i5 (.D(next_data_tx_7__N_378[5]), .CK(sys_clk), .CD(n52212), 
            .Q(data_tx[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam data_tx__i5.GSR = "ENABLED";
    FD1S3IX data_tx__i6 (.D(next_data_tx_7__N_378[6]), .CK(sys_clk), .CD(n52212), 
            .Q(data_tx[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam data_tx__i6.GSR = "ENABLED";
    FD1S3IX data_tx__i7 (.D(next_data_tx_7__N_378[7]), .CK(sys_clk), .CD(n52212), 
            .Q(data_tx[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam data_tx__i7.GSR = "ENABLED";
    LUT4 i26053_2_lut (.A(data_tx[2]), .B(\next_i2c_device_driver_state[0] ), 
         .Z(n19)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam i26053_2_lut.init = 16'h8888;
    LUT4 count_ms_15__I_0_875_i8_3_lut (.A(count_ms_15__N_910[4]), .B(count_ms_15__N_894[7]), 
         .C(n7654[7]), .Z(count_ms_15__N_396[7])) /* synthesis lut_function=(A (B (C))+!A (B+!(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(194[14] 219[12])
    defparam count_ms_15__I_0_875_i8_3_lut.init = 16'hc5c5;
    PFUMX i38678 (.BLUT(n22_adj_5328), .ALUT(n49472), .C0(n49693), .Z(next_data_tx_7__N_378[0]));
    PFUMX i38684 (.BLUT(n49477), .ALUT(n49478), .C0(\next_i2c_device_driver_state[4] ), 
          .Z(next_return_state_4__N_391[1]));
    PFUMX i67 (.BLUT(n48756), .ALUT(n48394), .C0(\i2c_top_debug[3] ), 
          .Z(n27_adj_5339));
    LUT4 count_ms_15__I_0_875_i7_3_lut (.A(count_ms_15__N_910[4]), .B(count_ms_15__N_894[6]), 
         .C(n7654[7]), .Z(count_ms_15__N_396[6])) /* synthesis lut_function=(A (B (C))+!A (B+!(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(194[14] 219[12])
    defparam count_ms_15__I_0_875_i7_3_lut.init = 16'hc5c5;
    PFUMX i62 (.BLUT(n24), .ALUT(n33), .C0(n49677), .Z(n36));
    PFUMX i40916 (.BLUT(n52483), .ALUT(n52484), .C0(\next_i2c_device_driver_return_state[1] ), 
          .Z(n52485));
    LUT4 i1_4_lut_adj_398 (.A(n34), .B(VL53L1X_measurement_period[5]), .C(VL53L1X_measurement_period[13]), 
         .D(measurement_period_tx_index[0]), .Z(n20)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_398.init = 16'ha088;
    LUT4 i25749_2_lut (.A(data_tx[5]), .B(\next_i2c_device_driver_state[0] ), 
         .Z(n19_adj_5268)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam i25749_2_lut.init = 16'h8888;
    PFUMX i40988 (.BLUT(n52591), .ALUT(n52592), .C0(data_reg[8]), .Z(n52593));
    LUT4 n33854_bdd_4_lut_40795_4_lut (.A(\next_i2c_device_driver_state[4] ), 
         .B(\next_i2c_device_driver_state[0] ), .C(n52201), .D(n33854), 
         .Z(n51719)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam n33854_bdd_4_lut_40795_4_lut.init = 16'h7340;
    LUT4 i1_4_lut_4_lut_adj_399 (.A(\next_i2c_device_driver_state[4] ), .B(\next_i2c_device_driver_state[3] ), 
         .C(n52440), .D(n7_adj_5301), .Z(n7240)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam i1_4_lut_4_lut_adj_399.init = 16'h5140;
    LUT4 i39207_3_lut_3_lut (.A(\next_i2c_device_driver_state[4] ), .B(n52157), 
         .C(n29_adj_5261), .Z(n49472)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam i39207_3_lut_3_lut.init = 16'he4e4;
    LUT4 i39136_3_lut (.A(n49495), .B(n52138), .C(\next_i2c_device_driver_state[3] ), 
         .Z(n49497)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam i39136_3_lut.init = 16'hcaca;
    CCU2D sub_257_add_2_5 (.A0(master_trigger_count_ms[3]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(master_trigger_count_ms[4]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n43797), .COUT(n43798), 
          .S0(n611[3]), .S1(n611[4]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(279[40:72])
    defparam sub_257_add_2_5.INIT0 = 16'h5555;
    defparam sub_257_add_2_5.INIT1 = 16'h5555;
    defparam sub_257_add_2_5.INJECT1_0 = "NO";
    defparam sub_257_add_2_5.INJECT1_1 = "NO";
    LUT4 i1_2_lut_2_lut_adj_400 (.A(\next_i2c_device_driver_state[4] ), .B(cal_reg_addr[0]), 
         .Z(n5_adj_5332)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam i1_2_lut_2_lut_adj_400.init = 16'h4444;
    LUT4 i19691_3_lut_rep_438 (.A(n30362), .B(n30361), .C(n30360), .Z(n52374)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19691_3_lut_rep_438.init = 16'hcaca;
    L6MUX21 i40090 (.D0(n50879), .D1(n50876), .SD(\next_i2c_device_driver_state[3] ), 
            .Z(next_target_read_count_5__N_414[1]));
    PFUMX i40088 (.BLUT(n50878), .ALUT(n50877), .C0(\next_i2c_device_driver_state[4] ), 
          .Z(n50879));
    LUT4 i1_2_lut_4_lut_adj_401 (.A(n30362), .B(n30361), .C(n30360), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_7__0__N_516)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_401.init = 16'hca00;
    LUT4 mux_3489_i2_3_lut_4_lut (.A(resetn_imu_N_1182), .B(next_addr_7__N_1168), 
         .C(n6974), .D(n6915[1]), .Z(next_VL53L1X_data_rx_reg_index[1])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(371[14:35])
    defparam mux_3489_i2_3_lut_4_lut.init = 16'h8f80;
    LUT4 mux_3489_i3_3_lut_4_lut (.A(resetn_imu_N_1182), .B(next_addr_7__N_1168), 
         .C(n6974), .D(n6915[2]), .Z(next_VL53L1X_data_rx_reg_index[2])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(371[14:35])
    defparam mux_3489_i3_3_lut_4_lut.init = 16'h8f80;
    LUT4 i2_3_lut_4_lut_adj_402 (.A(resetn_imu_N_1182), .B(next_addr_7__N_1168), 
         .C(n48249), .D(n52410), .Z(n53)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(371[14:35])
    defparam i2_3_lut_4_lut_adj_402.init = 16'h8000;
    CCU2D sub_257_add_2_3 (.A0(master_trigger_count_ms[1]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(master_trigger_count_ms[2]), 
          .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n43796), .COUT(n43797), 
          .S0(n611[1]), .S1(n611[2]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(279[40:72])
    defparam sub_257_add_2_3.INIT0 = 16'h5555;
    defparam sub_257_add_2_3.INIT1 = 16'h5555;
    defparam sub_257_add_2_3.INJECT1_0 = "NO";
    defparam sub_257_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_257_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(master_trigger_count_ms[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n43796), .S1(n611[0]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(279[40:72])
    defparam sub_257_add_2_1.INIT0 = 16'hF000;
    defparam sub_257_add_2_1.INIT1 = 16'h5555;
    defparam sub_257_add_2_1.INJECT1_0 = "NO";
    defparam sub_257_add_2_1.INJECT1_1 = "NO";
    PFUMX i40085 (.BLUT(n14_adj_5314), .ALUT(n50875), .C0(\next_i2c_device_driver_state[4] ), 
          .Z(n50876));
    CCU2D add_3739_17 (.A0(count_sys_clk_for_ms[15]), .B0(n14126), .C0(GND_net), 
          .D0(GND_net), .A1(count_sys_clk_for_ms[16]), .B1(count_ms[15]), 
          .C1(GND_net), .D1(GND_net), .CIN(n43794), .S0(count_sys_clk_for_ms_16__N_874[15]), 
          .S1(count_sys_clk_for_ms_16__N_874[16]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(211[14] 219[12])
    defparam add_3739_17.INIT0 = 16'h4444;
    defparam add_3739_17.INIT1 = 16'h7777;
    defparam add_3739_17.INJECT1_0 = "NO";
    defparam add_3739_17.INJECT1_1 = "NO";
    L6MUX21 i38621 (.D0(n49414), .D1(n49415), .SD(\next_i2c_device_driver_state[4] ), 
            .Z(next_data_reg_15__N_362[5]));
    LUT4 i1_2_lut_rep_524 (.A(\next_i2c_device_driver_state[4] ), .B(\next_i2c_device_driver_state[3] ), 
         .Z(n52460)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam i1_2_lut_rep_524.init = 16'h8888;
    CCU2D add_3739_15 (.A0(count_sys_clk_for_ms[13]), .B0(n14126), .C0(GND_net), 
          .D0(GND_net), .A1(count_sys_clk_for_ms[14]), .B1(n14126), .C1(GND_net), 
          .D1(GND_net), .CIN(n43793), .COUT(n43794), .S0(count_sys_clk_for_ms_16__N_874[13]), 
          .S1(count_sys_clk_for_ms_16__N_874[14]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(211[14] 219[12])
    defparam add_3739_15.INIT0 = 16'h7777;
    defparam add_3739_15.INIT1 = 16'h7777;
    defparam add_3739_15.INJECT1_0 = "NO";
    defparam add_3739_15.INJECT1_1 = "NO";
    PFUMX i40944 (.BLUT(n52525), .ALUT(n52526), .C0(\next_i2c_device_driver_state[2] ), 
          .Z(n24_adj_5322));
    LUT4 i27014_4_lut (.A(\next_data_tx_7__N_1032[1] ), .B(n37517), .C(data_tx[1]), 
         .D(\next_i2c_device_driver_state[0] ), .Z(n14_adj_5335)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(420[13] 870[20])
    defparam i27014_4_lut.init = 16'hc088;
    LUT4 i1_2_lut_3_lut_4_lut_adj_403 (.A(\next_i2c_device_driver_state[4] ), 
         .B(\next_i2c_device_driver_state[3] ), .C(\next_i2c_device_driver_state[0] ), 
         .D(n53892), .Z(n76)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam i1_2_lut_3_lut_4_lut_adj_403.init = 16'h0080;
    LUT4 count_ms_15__I_0_875_i10_3_lut (.A(count_ms_15__N_910[4]), .B(count_ms_15__N_894[9]), 
         .C(n7654[7]), .Z(count_ms_15__N_396[9])) /* synthesis lut_function=(A (B (C))+!A (B+!(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(194[14] 219[12])
    defparam count_ms_15__I_0_875_i10_3_lut.init = 16'hc5c5;
    LUT4 i2_2_lut_rep_367_3_lut (.A(\next_i2c_device_driver_state[4] ), .B(\next_i2c_device_driver_state[3] ), 
         .C(\next_i2c_device_driver_state[2] ), .Z(n52303)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam i2_2_lut_rep_367_3_lut.init = 16'h8080;
    LUT4 i2_2_lut_3_lut_4_lut (.A(\next_i2c_device_driver_state[4] ), .B(\next_i2c_device_driver_state[3] ), 
         .C(read_write_in), .D(\next_i2c_device_driver_state[2] ), .Z(n7_adj_5271)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam i2_2_lut_3_lut_4_lut.init = 16'h0800;
    L6MUX21 i38675 (.D0(n49468), .D1(n49469), .SD(\next_i2c_device_driver_state[4] ), 
            .Z(next_return_state_4__N_391[3]));
    LUT4 i19687_3_lut_rep_440 (.A(n30358), .B(n30357), .C(n30356), .Z(n52376)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i19687_3_lut_rep_440.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_404 (.A(n30358), .B(n30357), .C(n30356), .D(n52412), 
         .Z(VL53L1X_data_rx_reg_7__1__N_510)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam i1_2_lut_4_lut_adj_404.init = 16'hca00;
    LUT4 i1_2_lut_rep_529 (.A(resetn), .B(wd_event_active), .Z(next_addr_7__N_1168)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(371[14:35])
    defparam i1_2_lut_rep_529.init = 16'h2222;
    FD1P3JX master_trigger_count_ms_i6 (.D(master_trigger_count_ms_20__N_997[6]), 
            .SP(sys_clk_enable_224), .PD(n52182), .CK(sys_clk), .Q(master_trigger_count_ms[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(268[14] 281[12])
    defparam master_trigger_count_ms_i6.GSR = "ENABLED";
    FD1S3IX delay_timer_at_init_489 (.D(n48986), .CK(sys_clk_N_413), .CD(\next_i2c_device_driver_state[1] ), 
            .Q(delay_timer_at_init)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam delay_timer_at_init_489.GSR = "ENABLED";
    FD1P3JX master_trigger_count_ms_i7 (.D(master_trigger_count_ms_20__N_997[7]), 
            .SP(sys_clk_enable_224), .PD(n52182), .CK(sys_clk), .Q(master_trigger_count_ms[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(268[14] 281[12])
    defparam master_trigger_count_ms_i7.GSR = "ENABLED";
    FD1P3JX master_trigger_count_ms_i11 (.D(master_trigger_count_ms_20__N_997[11]), 
            .SP(sys_clk_enable_224), .PD(n52182), .CK(sys_clk), .Q(master_trigger_count_ms[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(268[14] 281[12])
    defparam master_trigger_count_ms_i11.GSR = "ENABLED";
    FD1P3JX master_trigger_count_ms_i12 (.D(master_trigger_count_ms_20__N_997[12]), 
            .SP(sys_clk_enable_224), .PD(n52182), .CK(sys_clk), .Q(master_trigger_count_ms[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(268[14] 281[12])
    defparam master_trigger_count_ms_i12.GSR = "ENABLED";
    FD1P3JX master_trigger_count_ms_i15 (.D(master_trigger_count_ms_20__N_997[15]), 
            .SP(sys_clk_enable_224), .PD(n52182), .CK(sys_clk), .Q(master_trigger_count_ms[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(268[14] 281[12])
    defparam master_trigger_count_ms_i15.GSR = "ENABLED";
    FD1P3JX master_trigger_count_ms_i16 (.D(master_trigger_count_ms_20__N_997[16]), 
            .SP(sys_clk_enable_224), .PD(n52182), .CK(sys_clk), .Q(master_trigger_count_ms[16])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(268[14] 281[12])
    defparam master_trigger_count_ms_i16.GSR = "ENABLED";
    FD1P3JX master_trigger_count_ms_i17 (.D(master_trigger_count_ms_20__N_997[17]), 
            .SP(sys_clk_enable_224), .PD(n52182), .CK(sys_clk), .Q(master_trigger_count_ms[17])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(268[14] 281[12])
    defparam master_trigger_count_ms_i17.GSR = "ENABLED";
    FD1P3JX master_trigger_count_ms_i19 (.D(master_trigger_count_ms_20__N_997[19]), 
            .SP(sys_clk_enable_224), .PD(n52182), .CK(sys_clk), .Q(master_trigger_count_ms[19])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(268[14] 281[12])
    defparam master_trigger_count_ms_i19.GSR = "ENABLED";
    PFUMX i40477 (.BLUT(n51507), .ALUT(n51506), .C0(measurement_period_tx_index[0]), 
          .Z(n51508));
    CCU2D add_3739_13 (.A0(count_sys_clk_for_ms[11]), .B0(n14126), .C0(GND_net), 
          .D0(GND_net), .A1(count_sys_clk_for_ms[12]), .B1(n14126), .C1(GND_net), 
          .D1(GND_net), .CIN(n43792), .COUT(n43793), .S0(count_sys_clk_for_ms_16__N_874[11]), 
          .S1(count_sys_clk_for_ms_16__N_874[12]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(211[14] 219[12])
    defparam add_3739_13.INIT0 = 16'h7777;
    defparam add_3739_13.INIT1 = 16'h4444;
    defparam add_3739_13.INJECT1_0 = "NO";
    defparam add_3739_13.INJECT1_1 = "NO";
    FD1S3IX delay_timer_done_487 (.D(n21625), .CK(sys_clk_N_413), .CD(n30677), 
            .Q(next_i2c_state_4__N_1050[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(174[14] 219[12])
    defparam delay_timer_done_487.GSR = "ENABLED";
    FD1P3AX measurement_period_tx_index_i1 (.D(next_measurement_period_tx_index[1]), 
            .SP(sys_clk_enable_242), .CK(sys_clk), .Q(measurement_period_tx_index[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam measurement_period_tx_index_i1.GSR = "ENABLED";
    FD1P3IX rx_from_VL53L1X_738 (.D(n13181[1]), .SP(sys_clk_enable_254), 
            .CD(n53891), .CK(sys_clk), .Q(rx_from_VL53L1X)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam rx_from_VL53L1X_738.GSR = "ENABLED";
    FD1P3AX measurement_period_tx_index_i0 (.D(next_measurement_period_tx_index[0]), 
            .SP(sys_clk_enable_255), .CK(sys_clk), .Q(measurement_period_tx_index[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam measurement_period_tx_index_i0.GSR = "ENABLED";
    FD1P3AX target_read_count_i0 (.D(next_target_read_count[0]), .SP(sys_clk_enable_256), 
            .CK(sys_clk), .Q(target_read_count[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam target_read_count_i0.GSR = "ENABLED";
    FD1S3IX go_730 (.D(n49101), .CK(sys_clk), .CD(n52421), .Q(go)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(347[14] 365[12])
    defparam go_730.GSR = "ENABLED";
    FD1S3AX valid_strobe_721 (.D(valid_strobe_N_1132), .CK(sys_clk), .Q(next_imu_data_valid)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(291[14] 304[12])
    defparam valid_strobe_721.GSR = "ENABLED";
    FD1S3DX VL53L1X_data_rx_reg_index_i0_i1_19946_19947_reset (.D(n23[1]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_index_5__N_460), .Q(n30619)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(229[14] 230[75])
    defparam VL53L1X_data_rx_reg_index_i0_i1_19946_19947_reset.GSR = "DISABLED";
    FD1S3BX VL53L1X_data_rx_reg_index_i0_i1_19946_19947_set (.D(n23[1]), .CK(sys_clk), 
            .PD(VL53L1X_data_rx_reg_index_5__N_442), .Q(n30618)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(229[14] 230[75])
    defparam VL53L1X_data_rx_reg_index_i0_i1_19946_19947_set.GSR = "DISABLED";
    FD1S3DX VL53L1X_data_rx_reg_index_i0_i2_19942_19943_reset (.D(n23[2]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_index_5__N_457), .Q(n30615)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(229[14] 230[75])
    defparam VL53L1X_data_rx_reg_index_i0_i2_19942_19943_reset.GSR = "DISABLED";
    FD1S3BX VL53L1X_data_rx_reg_index_i0_i2_19942_19943_set (.D(n23[2]), .CK(sys_clk), 
            .PD(VL53L1X_data_rx_reg_index_5__N_439), .Q(n30614)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(229[14] 230[75])
    defparam VL53L1X_data_rx_reg_index_i0_i2_19942_19943_set.GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_0[[0__718_19849_19850_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[0]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_0__0__N_774), .Q(n30522)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_0[[0__718_19849_19850_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_0[[0__718_19849_19850_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[0]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_0__0__N_772), .Q(n30521)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_0[[0__718_19849_19850_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_0[[1__714_19845_19846_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[1]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_0__1__N_768), .Q(n30518)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_0[[1__714_19845_19846_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_0[[1__714_19845_19846_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[1]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_0__1__N_766), .Q(n30517)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_0[[1__714_19845_19846_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_0[[2__710_19841_19842_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[2]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_0__2__N_762), .Q(n30514)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_0[[2__710_19841_19842_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_0[[2__710_19841_19842_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[2]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_0__2__N_760), .Q(n30513)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_0[[2__710_19841_19842_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_0[[3__706_19837_19838_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[3]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_0__3__N_756), .Q(n30510)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_0[[3__706_19837_19838_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_0[[3__706_19837_19838_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[3]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_0__3__N_754), .Q(n30509)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_0[[3__706_19837_19838_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_0[[4__702_19833_19834_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[4]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_0__4__N_750), .Q(n30506)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_0[[4__702_19833_19834_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_0[[4__702_19833_19834_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[4]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_0__4__N_748), .Q(n30505)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_0[[4__702_19833_19834_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_0[[5__698_19829_19830_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[5]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_0__5__N_744), .Q(n30502)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_0[[5__698_19829_19830_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_0[[5__698_19829_19830_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[5]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_0__5__N_742), .Q(n30501)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_0[[5__698_19829_19830_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_0[[6__694_19825_19826_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[6]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_0__6__N_738), .Q(n30498)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_0[[6__694_19825_19826_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_0[[6__694_19825_19826_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[6]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_0__6__N_736), .Q(n30497)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_0[[6__694_19825_19826_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_0[[7__690_19821_19822_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[7]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_0__7__N_732), .Q(n30494)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_0[[7__690_19821_19822_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_0[[7__690_19821_19822_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[7]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_0__7__N_730), .Q(n30493)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_0[[7__690_19821_19822_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_1[[0__686_19817_19818_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[8]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_1__0__N_726), .Q(n30490)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_1[[0__686_19817_19818_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_1[[0__686_19817_19818_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[8]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_1__0__N_724), .Q(n30489)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_1[[0__686_19817_19818_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_1[[1__682_19813_19814_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[9]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_1__1__N_720), .Q(n30486)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_1[[1__682_19813_19814_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_1[[1__682_19813_19814_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[9]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_1__1__N_718), .Q(n30485)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_1[[1__682_19813_19814_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_1[[2__678_19809_19810_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[10]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_1__2__N_714), .Q(n30482)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_1[[2__678_19809_19810_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_1[[2__678_19809_19810_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[10]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_1__2__N_712), .Q(n30481)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_1[[2__678_19809_19810_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_1[[3__674_19805_19806_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[11]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_1__3__N_708), .Q(n30478)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_1[[3__674_19805_19806_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_1[[3__674_19805_19806_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[11]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_1__3__N_706), .Q(n30477)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_1[[3__674_19805_19806_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_1[[4__670_19801_19802_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[12]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_1__4__N_702), .Q(n30474)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_1[[4__670_19801_19802_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_1[[4__670_19801_19802_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[12]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_1__4__N_700), .Q(n30473)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_1[[4__670_19801_19802_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_1[[5__666_19797_19798_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[13]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_1__5__N_696), .Q(n30470)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_1[[5__666_19797_19798_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_1[[5__666_19797_19798_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[13]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_1__5__N_694), .Q(n30469)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_1[[5__666_19797_19798_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_1[[6__662_19793_19794_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[14]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_1__6__N_690), .Q(n30466)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_1[[6__662_19793_19794_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_1[[6__662_19793_19794_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[14]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_1__6__N_688), .Q(n30465)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_1[[6__662_19793_19794_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_1[[7__658_19789_19790_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[15]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_1__7__N_684), .Q(n30462)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_1[[7__658_19789_19790_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_1[[7__658_19789_19790_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[15]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_1__7__N_682), .Q(n30461)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_1[[7__658_19789_19790_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_4[[0__638_19785_19786_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[32]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_4__0__N_662), .Q(n30458)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_4[[0__638_19785_19786_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_4[[0__638_19785_19786_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[32]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_4__0__N_660), .Q(n30457)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_4[[0__638_19785_19786_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_4[[1__634_19781_19782_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[33]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_4__1__N_656), .Q(n30454)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_4[[1__634_19781_19782_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_4[[1__634_19781_19782_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[33]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_4__1__N_654), .Q(n30453)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_4[[1__634_19781_19782_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_4[[2__630_19777_19778_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[34]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_4__2__N_650), .Q(n30450)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_4[[2__630_19777_19778_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_4[[2__630_19777_19778_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[34]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_4__2__N_648), .Q(n30449)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_4[[2__630_19777_19778_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_4[[3__626_19773_19774_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[35]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_4__3__N_644), .Q(n30446)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_4[[3__626_19773_19774_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_4[[3__626_19773_19774_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[35]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_4__3__N_642), .Q(n30445)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_4[[3__626_19773_19774_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_4[[4__622_19769_19770_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[36]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_4__4__N_638), .Q(n30442)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_4[[4__622_19769_19770_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_4[[4__622_19769_19770_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[36]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_4__4__N_636), .Q(n30441)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_4[[4__622_19769_19770_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_4[[5__618_19765_19766_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[37]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_4__5__N_632), .Q(n30438)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_4[[5__618_19765_19766_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_4[[5__618_19765_19766_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[37]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_4__5__N_630), .Q(n30437)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_4[[5__618_19765_19766_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_4[[6__614_19761_19762_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[38]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_4__6__N_626), .Q(n30434)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_4[[6__614_19761_19762_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_4[[6__614_19761_19762_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[38]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_4__6__N_624), .Q(n30433)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_4[[6__614_19761_19762_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_4[[7__610_19757_19758_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[39]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_4__7__N_620), .Q(n30430)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_4[[7__610_19757_19758_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_4[[7__610_19757_19758_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[39]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_4__7__N_618), .Q(n30429)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_4[[7__610_19757_19758_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_5[[0__606_19753_19754_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[40]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_5__0__N_614), .Q(n30426)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_5[[0__606_19753_19754_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_5[[0__606_19753_19754_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[40]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_5__0__N_612), .Q(n30425)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_5[[0__606_19753_19754_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_5[[1__602_19749_19750_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[41]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_5__1__N_608), .Q(n30422)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_5[[1__602_19749_19750_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_5[[1__602_19749_19750_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[41]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_5__1__N_606), .Q(n30421)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_5[[1__602_19749_19750_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_5[[2__598_19745_19746_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[42]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_5__2__N_602), .Q(n30418)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_5[[2__598_19745_19746_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_5[[2__598_19745_19746_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[42]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_5__2__N_600), .Q(n30417)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_5[[2__598_19745_19746_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_5[[3__594_19741_19742_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[43]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_5__3__N_596), .Q(n30414)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_5[[3__594_19741_19742_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_5[[3__594_19741_19742_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[43]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_5__3__N_594), .Q(n30413)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_5[[3__594_19741_19742_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_5[[4__590_19737_19738_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[44]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_5__4__N_590), .Q(n30410)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_5[[4__590_19737_19738_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_5[[4__590_19737_19738_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[44]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_5__4__N_588), .Q(n30409)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_5[[4__590_19737_19738_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_5[[5__586_19733_19734_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[45]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_5__5__N_584), .Q(n30406)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_5[[5__586_19733_19734_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_5[[5__586_19733_19734_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[45]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_5__5__N_582), .Q(n30405)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_5[[5__586_19733_19734_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_5[[6__582_19729_19730_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[46]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_5__6__N_578), .Q(n30402)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_5[[6__582_19729_19730_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_5[[6__582_19729_19730_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[46]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_5__6__N_576), .Q(n30401)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_5[[6__582_19729_19730_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_5[[7__578_19725_19726_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[47]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_5__7__N_572), .Q(n30398)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_5[[7__578_19725_19726_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_5[[7__578_19725_19726_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[47]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_5__7__N_570), .Q(n30397)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_5[[7__578_19725_19726_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_6[[0__574_19721_19722_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[48]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_6__0__N_566), .Q(n30394)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_6[[0__574_19721_19722_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_6[[0__574_19721_19722_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[48]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_6__0__N_564), .Q(n30393)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_6[[0__574_19721_19722_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_6[[1__570_19717_19718_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[49]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_6__1__N_560), .Q(n30390)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_6[[1__570_19717_19718_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_6[[1__570_19717_19718_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[49]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_6__1__N_558), .Q(n30389)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_6[[1__570_19717_19718_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_6[[2__566_19713_19714_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[50]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_6__2__N_554), .Q(n30386)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_6[[2__566_19713_19714_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_6[[2__566_19713_19714_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[50]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_6__2__N_552), .Q(n30385)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_6[[2__566_19713_19714_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_6[[3__562_19709_19710_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[51]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_6__3__N_548), .Q(n30382)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_6[[3__562_19709_19710_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_6[[3__562_19709_19710_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[51]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_6__3__N_546), .Q(n30381)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_6[[3__562_19709_19710_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_6[[4__558_19705_19706_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[52]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_6__4__N_542), .Q(n30378)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_6[[4__558_19705_19706_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_6[[4__558_19705_19706_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[52]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_6__4__N_540), .Q(n30377)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_6[[4__558_19705_19706_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_6[[5__554_19701_19702_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[53]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_6__5__N_536), .Q(n30374)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_6[[5__554_19701_19702_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_6[[5__554_19701_19702_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[53]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_6__5__N_534), .Q(n30373)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_6[[5__554_19701_19702_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_6[[6__550_19697_19698_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[54]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_6__6__N_530), .Q(n30370)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_6[[6__550_19697_19698_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_6[[6__550_19697_19698_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[54]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_6__6__N_528), .Q(n30369)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_6[[6__550_19697_19698_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_6[[7__546_19693_19694_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[55]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_6__7__N_524), .Q(n30366)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_6[[7__546_19693_19694_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_6[[7__546_19693_19694_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[55]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_6__7__N_522), .Q(n30365)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_6[[7__546_19693_19694_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_7[[0__542_19689_19690_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[56]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_7__0__N_518), .Q(n30362)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_7[[0__542_19689_19690_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_7[[0__542_19689_19690_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[56]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_7__0__N_516), .Q(n30361)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_7[[0__542_19689_19690_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_7[[1__538_19685_19686_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[57]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_7__1__N_512), .Q(n30358)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_7[[1__538_19685_19686_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_7[[1__538_19685_19686_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[57]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_7__1__N_510), .Q(n30357)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_7[[1__538_19685_19686_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_7[[2__534_19681_19682_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[58]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_7__2__N_506), .Q(n30354)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_7[[2__534_19681_19682_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_7[[2__534_19681_19682_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[58]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_7__2__N_504), .Q(n30353)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_7[[2__534_19681_19682_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_7[[3__530_19677_19678_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[59]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_7__3__N_500), .Q(n30350)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_7[[3__530_19677_19678_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_7[[3__530_19677_19678_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[59]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_7__3__N_498), .Q(n30349)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_7[[3__530_19677_19678_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_7[[4__526_19673_19674_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[60]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_7__4__N_494), .Q(n30346)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_7[[4__526_19673_19674_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_7[[4__526_19673_19674_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[60]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_7__4__N_492), .Q(n30345)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_7[[4__526_19673_19674_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_7[[5__522_19669_19670_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[61]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_7__5__N_488), .Q(n30342)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_7[[5__522_19669_19670_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_7[[5__522_19669_19670_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[61]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_7__5__N_486), .Q(n30341)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_7[[5__522_19669_19670_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_7[[6__518_19665_19666_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[62]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_7__6__N_482), .Q(n30338)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_7[[6__518_19665_19666_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_7[[6__518_19665_19666_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[62]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_7__6__N_480), .Q(n30337)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_7[[6__518_19665_19666_set .GSR = "DISABLED";
    FD1S3DX \VL53L1X_data_rx_reg_7[[7__514_19661_19662_reset  (.D(VL53L1X_data_rx_reg_7__7__N_472[63]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_7__7__N_476), .Q(n30334)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_7[[7__514_19661_19662_reset .GSR = "DISABLED";
    FD1S3BX \VL53L1X_data_rx_reg_7[[7__514_19661_19662_set  (.D(VL53L1X_data_rx_reg_7__7__N_472[63]), 
            .CK(sys_clk), .PD(VL53L1X_data_rx_reg_7__7__N_473), .Q(n30333)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(251[14] 253[12])
    defparam \VL53L1X_data_rx_reg_7[[7__514_19661_19662_set .GSR = "DISABLED";
    FD1S3DX VL53L1X_data_rx_reg_index_i0_i0_19657_19658_reset (.D(n23[0]), 
            .CK(sys_clk), .CD(VL53L1X_data_rx_reg_index_5__N_463), .Q(n30330)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(229[14] 230[75])
    defparam VL53L1X_data_rx_reg_index_i0_i0_19657_19658_reset.GSR = "DISABLED";
    FD1S3BX VL53L1X_data_rx_reg_index_i0_i0_19657_19658_set (.D(n23[0]), .CK(sys_clk), 
            .PD(VL53L1X_data_rx_reg_index_5__N_445), .Q(n30329)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=9, LSE_RCOL=6, LSE_LLINE=299, LSE_RLINE=349 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(229[14] 230[75])
    defparam VL53L1X_data_rx_reg_index_i0_i0_19657_19658_set.GSR = "DISABLED";
    FD1S1D i19656 (.D(n53885), .CK(VL53L1X_data_rx_reg_index_5__N_445), 
           .CD(VL53L1X_data_rx_reg_index_5__N_463), .Q(n30328));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(229[14] 230[75])
    defparam i19656.GSR = "DISABLED";
    i2c_module i2c (.\i2c_top_debug[0] (\i2c_top_debug[0] ), .\i2c_top_debug[1] (\i2c_top_debug[1] ), 
            .n53886(n53886), .\i2c_top_debug[2] (i2c_top_debug[2]), .\i2c_top_debug[3] (\i2c_top_debug[3] ), 
            .\i2c_top_debug[4] (\i2c_top_debug[4] ), .n53892(n53892), .\next_i2c_device_driver_state[0] (\next_i2c_device_driver_state[0] ), 
            .\next_i2c_device_driver_state[2] (\next_i2c_device_driver_state[2] ), 
            .\data_reg[5] (data_reg[5]), .n29(n29_adj_5298), .n52425(n52425), 
            .\i2c_top_debug[5] (\i2c_top_debug[5] ), .resetn_derived_2(resetn_derived_2), 
            .n53885(n53885), .sys_clk(sys_clk), .wd_event_active(wd_event_active), 
            .data_rx({data_rx}), .\data_reg[7] (data_reg[7]), .n27301(n27301), 
            .one_byte_ready(one_byte_ready), .next_addr_7__N_1168(next_addr_7__N_1168), 
            .read_write_in(read_write_in), .byte_rd_left_5__N_1255(byte_rd_left_5__N_1255), 
            .n52142(n52142), .n45689(n45689), .resetn_imu_N_1182(resetn_imu_N_1182), 
            .n6(n6_adj_5333), .\next_i2c_device_driver_state[3] (\next_i2c_device_driver_state[3] ), 
            .n46519(n46519), .n46521(n46521), .n52205(n52205), .n52306(n52306), 
            .n66(n66), .n52318(n52318), .n52188(n52188), .\data_reg[1] (data_reg[1]), 
            .n10(n10_adj_5276), .is_2_byte_reg(is_2_byte_reg), .\target_read_count[0] (target_read_count[0]), 
            .\data_reg[2] (data_reg[2]), .data_tx({data_tx}), .n51003(n51003), 
            .n27391(n27391), .\data_reg[3] (data_reg[3]), .\data_reg[4] (data_reg[4]), 
            .\target_read_count[1] (target_read_count[1]), .n48722(n48722), 
            .n48394(n48394), .n52248(n52248), .n47760(n47760), .\next_i2c_state_4__N_1050[0] (next_i2c_state_4__N_1050[0]), 
            .n69(n69), .clear_waiting_ms_N_893(n2485[7]), .clear_waiting_ms(n7654[7]), 
            .\next_i2c_device_driver_state[4] (\next_i2c_device_driver_state[4] ), 
            .n7(n7_adj_5278), .n34018(n34018), .go(go), .GND_net(GND_net), 
            .n48829(n48829), .n33(n33), .\data_reg[6] (data_reg[6]), .n48756(n48756), 
            .n7246(n7246), .n49365(n49365), .resetn(resetn), .\data_reg[0] (data_reg[0]), 
            .n48496(n48496), .n52450(n52450), .delay_timer_at_init(delay_timer_at_init), 
            .\next_i2c_state_4__N_1090[0] (next_i2c_state_4__N_1090[0]), .n1(n1_adj_5338), 
            .n1_adj_1(n1_adj_5324), .\data_reg[8] (data_reg[8]), .n52140(n52140), 
            .\next_data_reg_15__N_362[0] (next_data_reg_15__N_362[0]), .n48098(n48098), 
            .i2c2_sdaoen(i2c2_sdaoen), .i2c2_sdao(i2c2_sdao), .i2c2_scloen(i2c2_scloen), 
            .i2c2_sclo(i2c2_sclo), .i2c2_sdai(i2c2_sdai), .i2c2_scli(i2c2_scli), 
            .i2c1_sdaoen(i2c1_sdaoen), .i2c1_sdao(i2c1_sdao), .i2c1_scloen(i2c1_scloen), 
            .i2c1_sclo(i2c1_sclo), .i2c1_sdai(i2c1_sdai), .i2c1_scli(i2c1_scli), 
            .VCC_net(VCC_net)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(140[16] 159[6])
    
endmodule
//
// Verilog Description of module i2c_module
//

module i2c_module (\i2c_top_debug[0] , \i2c_top_debug[1] , n53886, \i2c_top_debug[2] , 
            \i2c_top_debug[3] , \i2c_top_debug[4] , n53892, \next_i2c_device_driver_state[0] , 
            \next_i2c_device_driver_state[2] , \data_reg[5] , n29, n52425, 
            \i2c_top_debug[5] , resetn_derived_2, n53885, sys_clk, wd_event_active, 
            data_rx, \data_reg[7] , n27301, one_byte_ready, next_addr_7__N_1168, 
            read_write_in, byte_rd_left_5__N_1255, n52142, n45689, resetn_imu_N_1182, 
            n6, \next_i2c_device_driver_state[3] , n46519, n46521, n52205, 
            n52306, n66, n52318, n52188, \data_reg[1] , n10, is_2_byte_reg, 
            \target_read_count[0] , \data_reg[2] , data_tx, n51003, 
            n27391, \data_reg[3] , \data_reg[4] , \target_read_count[1] , 
            n48722, n48394, n52248, n47760, \next_i2c_state_4__N_1050[0] , 
            n69, clear_waiting_ms_N_893, clear_waiting_ms, \next_i2c_device_driver_state[4] , 
            n7, n34018, go, GND_net, n48829, n33, \data_reg[6] , 
            n48756, n7246, n49365, resetn, \data_reg[0] , n48496, 
            n52450, delay_timer_at_init, \next_i2c_state_4__N_1090[0] , 
            n1, n1_adj_1, \data_reg[8] , n52140, \next_data_reg_15__N_362[0] , 
            n48098, i2c2_sdaoen, i2c2_sdao, i2c2_scloen, i2c2_sclo, 
            i2c2_sdai, i2c2_scli, i2c1_sdaoen, i2c1_sdao, i2c1_scloen, 
            i2c1_sclo, i2c1_sdai, i2c1_scli, VCC_net) /* synthesis syn_module_defined=1 */ ;
    output \i2c_top_debug[0] ;
    output \i2c_top_debug[1] ;
    output n53886;
    output \i2c_top_debug[2] ;
    output \i2c_top_debug[3] ;
    output \i2c_top_debug[4] ;
    input n53892;
    input \next_i2c_device_driver_state[0] ;
    input \next_i2c_device_driver_state[2] ;
    input \data_reg[5] ;
    output n29;
    output n52425;
    output \i2c_top_debug[5] ;
    input resetn_derived_2;
    input n53885;
    input sys_clk;
    output wd_event_active;
    output [7:0]data_rx;
    input \data_reg[7] ;
    output n27301;
    output one_byte_ready;
    input next_addr_7__N_1168;
    input read_write_in;
    input byte_rd_left_5__N_1255;
    output n52142;
    input n45689;
    output resetn_imu_N_1182;
    input n6;
    input \next_i2c_device_driver_state[3] ;
    input n46519;
    input n46521;
    input n52205;
    output n52306;
    output n66;
    input n52318;
    output n52188;
    input \data_reg[1] ;
    input n10;
    input is_2_byte_reg;
    input \target_read_count[0] ;
    input \data_reg[2] ;
    input [7:0]data_tx;
    output n51003;
    input n27391;
    input \data_reg[3] ;
    input \data_reg[4] ;
    input \target_read_count[1] ;
    output n48722;
    output n48394;
    output n52248;
    input n47760;
    input \next_i2c_state_4__N_1050[0] ;
    output n69;
    input clear_waiting_ms_N_893;
    output clear_waiting_ms;
    input \next_i2c_device_driver_state[4] ;
    output n7;
    output n34018;
    input go;
    input GND_net;
    output n48829;
    output n33;
    input \data_reg[6] ;
    output n48756;
    input n7246;
    output n49365;
    input resetn;
    input \data_reg[0] ;
    input n48496;
    input n52450;
    input delay_timer_at_init;
    input \next_i2c_state_4__N_1090[0] ;
    output n1;
    output n1_adj_1;
    input \data_reg[8] ;
    input n52140;
    output \next_data_reg_15__N_362[0] ;
    input n48098;
    output i2c2_sdaoen;
    output i2c2_sdao;
    output i2c2_scloen;
    output i2c2_sclo;
    input i2c2_sdai;
    input i2c2_scli;
    output i2c1_sdaoen;
    output i2c1_sdao;
    output i2c1_scloen;
    output i2c1_sclo;
    input i2c1_sdai;
    input i2c1_scli;
    input VCC_net;
    
    wire sys_clk /* synthesis SET_AS_NETWORK=sys_clk, is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(220[10:17])
    wire next_addr_7__N_1168 /* synthesis is_clock=1, SET_AS_NETWORK=\I2C_Devices/i2c/next_addr_7__N_1168 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(45[15:24])
    wire data_latch /* synthesis is_clock=1, SET_AS_NETWORK=\I2C_Devices/i2c/data_latch */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(56[10:20])
    wire next_ack_flag_N_1498 /* synthesis is_clock=1, SET_AS_NETWORK=\I2C_Devices/i2c/next_ack_flag_N_1498 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(55[20:33])
    wire i2c2_scli /* synthesis is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_efb_wb.v(34[10:19])
    wire i2c1_scli /* synthesis is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_efb_wb.v(40[10:19])
    
    wire n26115, n48875, n48712, n76, n38227, n37916, n52432, 
        n38303, n52230, n4, n30, count_us_11__N_1299, n52424, n6_c, 
        n49387, n26272, n49767, n51038, n51035, n51040, n50987, 
        n49034, n28215, n51037, n26271, n52025, n30594, count_us_11__N_1215;
    wire [5:0]next_i2c_cmd_state_5__N_1479;
    
    wire n49519, n52608, n51536, n43987, n43988, n43989, n4068, 
        n52229, n4_adj_5200, n49417, n52538, n52537, module_data_out_7__N_1332;
    wire [7:0]data_rx_adj_5257;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(37[16:23])
    
    wire n51194, n10_c, n23, n24, n49498, n51036, n30621, byte_rd_left_5__N_1266, 
        byte_rd_left_5__N_1282, n48963, n29_adj_5202, n49391;
    wire [31:0]count_wd_delay;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(51[16:30])
    wire [31:0]count_wd_delay_31__N_1216;
    wire [7:0]addr;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(35[16:20])
    wire [7:0]next_addr;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(45[15:24])
    
    wire we, next_we, stb, next_stb;
    wire [7:0]data_tx_c;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(36[16:23])
    wire [7:0]next_data_tx;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(46[15:27])
    
    wire ack_flag, next_ack_flag, next_one_byte_ready, n31, read_action, 
        read_write_in_N_1023, write_action;
    wire [7:0]next_addr_7__N_1160;
    wire [5:0]byte_rd_left;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(58[15:27])
    wire [5:0]byte_rd_left_5__N_1248;
    
    wire n52287, n7628, n52175;
    wire [1:0]n12358;
    
    wire n30625, byte_rd_left_5__N_1265, byte_rd_left_5__N_1279, next_data_latch_N_1505, 
        n32, n52466, n52241, n4_adj_5203, n25, n53177, n53178, 
        n53882, n21941, n21, n49459, n52193, n63;
    wire [31:0]n77;
    
    wire n48117, n15, n49064, n30_adj_5204, n31_adj_5205, n30623, 
        n30622, n52439, n52286, n32988, n52607, n47361, n52606, 
        n15_adj_5206, n18960, n31_adj_5207, n53172, n53173, n53883, 
        n53171, n51768, n51856, n51924, n49440, n51741, n49392, 
        n52452, n10_adj_5208, n49402, n49403, n51918, n51917, n53875, 
        n52228, n51738, n51740, n53872, n4_adj_5210, n52289, n52288, 
        sys_clk_enable_231, n52174;
    wire [8:0]n2486;
    
    wire n52200, n51764, n14, n51767, n51766, n52239, n1516, n19779, 
        n38357, n49768, n10_adj_5212, n52464, n50986;
    wire [1:0]byte_wr_left;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(59[15:27])
    wire [1:0]n2;
    
    wire n48107, n48108, n29_adj_5214, n26203, n51853, n52263, n50, 
        n52293, n49388, n48025, n49, n62, n58, n50_adj_5215, n41, 
        n60, n54, n42, n52, n38, n56, n46;
    wire [7:0]n1296;
    
    wire n37968, n24_adj_5217, n25_adj_5218, n37653, n49419, n49395, 
        n51921, n10_adj_5219, n12, n46343, n30627, n30626, n28, 
        n27058, n48426, n51854, n52273, n51855, n49_adj_5220, n51739, 
        n51922, n51923, n9, n52459, n5, n52024, n48, n62_adj_5221, 
        n52234, n33015, n22, n52455, n49460, n49461, n52316, n51852, 
        n51759, n51737, n4_adj_5222, n49516, n49518, n8, n30598;
    wire [11:0]n26;
    
    wire n52299;
    wire [1:0]n12368;
    
    wire n8_adj_5228, n30601, n30604, n30607;
    wire [11:0]count_us;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(49[16:24])
    
    wire count_us_11__N_1209;
    wire [11:0]count_us_11__N_1287;
    
    wire n30610, n49529, n7_c, n4_adj_5238, n52298, n51765, data_rx_7__N_1159, 
        n7_adj_5239, n53881, n49650, n52232, n52192, n48815, n51734, 
        n51849, n37453, n7_adj_5241, n49517, n31_adj_5242, n52416, 
        n49652, n52262, ack, sys_clk_enable_148;
    wire [1:0]n17;
    
    wire n49672, n48845, n52301, n29_adj_5243, n52423, n52275, n49394, 
        n49501, n38161, n48814, n52436, n52277, n45033, n50985, 
        n52431, n49502, n28051, n49505, n49504, n7_adj_5245, n52026, 
        n8_adj_5246, n52259, n52300, n49418, n8_adj_5247, n49393, 
        n49506, n52028, n52027, n49389, n31_adj_5248, n52291, n48112, 
        n52539, n43947, n43946, n29_adj_5249, n44475, n14_adj_5251, 
        n51851, n53, n14_adj_5253, n32969, n43945, n49503, n43944, 
        n49222, n49216, n43943, n43942, n49212, n30599, n30611, 
        n30602, n30605, n30596, n30595, n30608, clear_waiting_us, 
        n49438, n49439, n6849, n49390, n43925, n43924, n43923, 
        n43922, n43921, n43920;
    wire [31:0]count_wd_delay_31__N_1300;
    
    wire n53175, n43919, n43918, n43917, n43916, n43915, n43914, 
        n43913, n43912, n43911, n43910, n53176, n8_adj_5256;
    
    LUT4 i15635_3_lut_3_lut (.A(\i2c_top_debug[0] ), .B(\i2c_top_debug[1] ), 
         .C(n53886), .Z(n26115)) /* synthesis lut_function=(A ((C)+!B)+!A !((C)+!B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i15635_3_lut_3_lut.init = 16'ha6a6;
    PFUMX i78 (.BLUT(n48875), .ALUT(n48712), .C0(\i2c_top_debug[0] ), 
          .Z(n76));
    PFUMX i2c_top_debug_5__I_0_767_Mux_0_i29 (.BLUT(n38227), .ALUT(n37916), 
          .C0(n52432), .Z(n38303)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;
    LUT4 i2c_top_debug_5__I_0_768_Mux_0_i30_4_lut (.A(\i2c_top_debug[2] ), 
         .B(n52230), .C(\i2c_top_debug[3] ), .D(n4), .Z(n30)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i2c_top_debug_5__I_0_768_Mux_0_i30_4_lut.init = 16'hcac0;
    LUT4 i39330_3_lut_4_lut (.A(count_us_11__N_1299), .B(n52424), .C(\i2c_top_debug[2] ), 
         .D(n6_c), .Z(n49387)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam i39330_3_lut_4_lut.init = 16'hf808;
    LUT4 i2_4_lut_4_lut_4_lut (.A(\i2c_top_debug[3] ), .B(\i2c_top_debug[2] ), 
         .C(\i2c_top_debug[1] ), .D(\i2c_top_debug[4] ), .Z(n48875)) /* synthesis lut_function=(A (B (C+(D))+!B (D))+!A (B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam i2_4_lut_4_lut_4_lut.init = 16'hffd4;
    LUT4 i24311_4_lut_4_lut (.A(n53892), .B(\next_i2c_device_driver_state[0] ), 
         .C(\next_i2c_device_driver_state[2] ), .D(\data_reg[5] ), .Z(n29)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(B ((D)+!C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i24311_4_lut_4_lut.init = 16'h6404;
    LUT4 i39161_1_lut_4_lut (.A(\i2c_top_debug[4] ), .B(n26272), .C(n52425), 
         .D(n38303), .Z(n49767)) /* synthesis lut_function=(!(A (D)+!A (B+(C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i39161_1_lut_4_lut.init = 16'h01ab;
    LUT4 n51039_bdd_2_lut_4_lut (.A(n51038), .B(n51035), .C(\i2c_top_debug[2] ), 
         .D(\i2c_top_debug[5] ), .Z(n51040)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam n51039_bdd_2_lut_4_lut.init = 16'hffca;
    LUT4 n45_bdd_4_lut_40490_4_lut (.A(\i2c_top_debug[0] ), .B(\i2c_top_debug[1] ), 
         .C(\i2c_top_debug[4] ), .D(\i2c_top_debug[3] ), .Z(n51035)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+(D)))+!A !(B (C (D)+!C !(D))+!B !(C+(D))))) */ ;
    defparam n45_bdd_4_lut_40490_4_lut.init = 16'h622d;
    LUT4 i39187_3_lut (.A(n50987), .B(n49034), .C(\i2c_top_debug[5] ), 
         .Z(n28215)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i39187_3_lut.init = 16'hcaca;
    LUT4 n45_bdd_3_lut_40491_4_lut_3_lut (.A(\i2c_top_debug[0] ), .B(\i2c_top_debug[1] ), 
         .C(\i2c_top_debug[3] ), .Z(n51037)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)+!B !(C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam n45_bdd_3_lut_40491_4_lut_3_lut.init = 16'h4949;
    LUT4 i15785_3_lut_4_lut_3_lut (.A(\i2c_top_debug[0] ), .B(\i2c_top_debug[1] ), 
         .C(\i2c_top_debug[2] ), .Z(n26271)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B (C)+!B !(C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i15785_3_lut_4_lut_3_lut.init = 16'h4949;
    LUT4 next_data_tx_7__N_1439_4__bdd_2_lut_40820_4_lut_4_lut (.A(\i2c_top_debug[0] ), 
         .B(\i2c_top_debug[1] ), .C(\i2c_top_debug[2] ), .D(n52425), .Z(n52025)) /* synthesis lut_function=(!(A (B (C+(D))+!B ((D)+!C))+!A (B (D)+!B (C+(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam next_data_tx_7__N_1439_4__bdd_2_lut_40820_4_lut_4_lut.init = 16'h006d;
    FD1S1D i19922 (.D(n53885), .CK(resetn_derived_2), .CD(count_us_11__N_1215), 
           .Q(n30594));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(128[14] 131[34])
    defparam i19922.GSR = "DISABLED";
    FD1S3IX i2c_cmd_state__i1 (.D(next_i2c_cmd_state_5__N_1479[0]), .CK(sys_clk), 
            .CD(wd_event_active), .Q(\i2c_top_debug[0] )) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam i2c_cmd_state__i1.GSR = "ENABLED";
    LUT4 n49519_bdd_3_lut_40882 (.A(n49519), .B(n52608), .C(n53886), .Z(n51536)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n49519_bdd_3_lut_40882.init = 16'hcaca;
    PFUMX i33213 (.BLUT(n43987), .ALUT(n43988), .C0(\i2c_top_debug[1] ), 
          .Z(n43989));
    LUT4 i38622_4_lut (.A(n4068), .B(n52229), .C(\i2c_top_debug[3] ), 
         .D(n4_adj_5200), .Z(n49417)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i38622_4_lut.init = 16'hcac0;
    LUT4 i26818_4_lut_4_lut_then_4_lut (.A(n52425), .B(\i2c_top_debug[2] ), 
         .C(\i2c_top_debug[1] ), .D(\i2c_top_debug[0] ), .Z(n52538)) /* synthesis lut_function=(!(A+(B (C (D)+!C !(D))+!B !(C+!(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i26818_4_lut_4_lut_then_4_lut.init = 16'h1451;
    LUT4 i26818_4_lut_4_lut_else_4_lut (.A(n52425), .B(\i2c_top_debug[2] ), 
         .C(\i2c_top_debug[1] ), .D(\i2c_top_debug[0] ), .Z(n52537)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i26818_4_lut_4_lut_else_4_lut.init = 16'h4000;
    FD1P3AX module_data_out_i0_i0 (.D(data_rx_adj_5257[0]), .SP(module_data_out_7__N_1332), 
            .CK(sys_clk), .Q(data_rx[0])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(209[14] 216[12])
    defparam module_data_out_i0_i0.GSR = "ENABLED";
    LUT4 i2c_top_debug_5__I_0_768_Mux_7_i10_4_lut (.A(n51194), .B(\data_reg[7] ), 
         .C(\i2c_top_debug[1] ), .D(n27301), .Z(n10_c)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i2c_top_debug_5__I_0_768_Mux_7_i10_4_lut.init = 16'hca0a;
    PFUMX i38703 (.BLUT(n23), .ALUT(n24), .C0(\i2c_top_debug[1] ), .Z(n49498));
    LUT4 n45_bdd_3_lut_40191_3_lut (.A(\i2c_top_debug[0] ), .B(\i2c_top_debug[1] ), 
         .C(\i2c_top_debug[3] ), .Z(n51036)) /* synthesis lut_function=(A (B (C))+!A !(B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam n45_bdd_3_lut_40191_3_lut.init = 16'h9595;
    FD1S1D i19949 (.D(n53885), .CK(byte_rd_left_5__N_1266), .CD(byte_rd_left_5__N_1282), 
           .Q(n30621));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(225[14] 227[12])
    defparam i19949.GSR = "DISABLED";
    PFUMX i38596 (.BLUT(n48963), .ALUT(n29_adj_5202), .C0(\i2c_top_debug[3] ), 
          .Z(n49391));
    FD1S3AY count_wd_delay_i0 (.D(count_wd_delay_31__N_1216[0]), .CK(sys_clk), 
            .Q(count_wd_delay[0])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[14] 151[12])
    defparam count_wd_delay_i0.GSR = "ENABLED";
    FD1S3AX addr_i1 (.D(next_addr[0]), .CK(sys_clk), .Q(addr[0])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam addr_i1.GSR = "ENABLED";
    FD1S3AX we_688 (.D(next_we), .CK(sys_clk), .Q(we)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam we_688.GSR = "ENABLED";
    FD1S3AX stb_689 (.D(next_stb), .CK(sys_clk), .Q(stb)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam stb_689.GSR = "ENABLED";
    FD1S3AX data_tx_i0 (.D(next_data_tx[0]), .CK(sys_clk), .Q(data_tx_c[0])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam data_tx_i0.GSR = "ENABLED";
    FD1S3AX ack_flag_693 (.D(next_ack_flag), .CK(sys_clk), .Q(ack_flag)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam ack_flag_693.GSR = "ENABLED";
    FD1S3AX one_byte_ready_695 (.D(next_one_byte_ready), .CK(sys_clk), .Q(one_byte_ready)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam one_byte_ready_695.GSR = "ENABLED";
    FD1S1I next_data_tx_7__I_0_i1 (.D(n31), .CK(next_addr_7__N_1168), .CD(\i2c_top_debug[5] ), 
           .Q(next_data_tx[0])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(231[5] 1039[8])
    defparam next_data_tx_7__I_0_i1.GSR = "DISABLED";
    FD1S3AX read_action_699 (.D(read_write_in_N_1023), .CK(sys_clk), .Q(read_action)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(190[14] 199[12])
    defparam read_action_699.GSR = "ENABLED";
    FD1S3AX write_action_700 (.D(read_write_in), .CK(sys_clk), .Q(write_action)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(190[14] 199[12])
    defparam write_action_700.GSR = "ENABLED";
    FD1S3AX next_one_byte_ready_702 (.D(module_data_out_7__N_1332), .CK(sys_clk), 
            .Q(next_one_byte_ready)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(209[14] 216[12])
    defparam next_one_byte_ready_702.GSR = "ENABLED";
    FD1S1A next_addr_7__I_0_i1 (.D(next_addr_7__N_1160[0]), .CK(next_addr_7__N_1168), 
           .Q(next_addr[0])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(231[5] 1039[8])
    defparam next_addr_7__I_0_i1.GSR = "DISABLED";
    FD1S3DX byte_rd_left_i5 (.D(byte_rd_left_5__N_1248[5]), .CK(data_latch), 
            .CD(byte_rd_left_5__N_1255), .Q(byte_rd_left[5])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(225[14] 227[12])
    defparam byte_rd_left_i5.GSR = "DISABLED";
    FD1S3DX byte_rd_left_i4 (.D(byte_rd_left_5__N_1248[4]), .CK(data_latch), 
            .CD(byte_rd_left_5__N_1255), .Q(byte_rd_left[4])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(225[14] 227[12])
    defparam byte_rd_left_i4.GSR = "DISABLED";
    FD1S3DX byte_rd_left_i3 (.D(n52287), .CK(data_latch), .CD(byte_rd_left_5__N_1255), 
            .Q(byte_rd_left[3])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(225[14] 227[12])
    defparam byte_rd_left_i3.GSR = "DISABLED";
    FD1S1A next_stb_I_0 (.D(next_addr_7__N_1160[6]), .CK(next_addr_7__N_1168), 
           .Q(next_stb)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(231[5] 1039[8])
    defparam next_stb_I_0.GSR = "DISABLED";
    LUT4 mux_4861_i1_4_lut_4_lut (.A(n52425), .B(data_latch), .C(n7628), 
         .D(n52175), .Z(n12358[0])) /* synthesis lut_function=(!(A (B (C)+!B (D))+!A ((C)+!B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(976[30:91])
    defparam mux_4861_i1_4_lut_4_lut.init = 16'h0c2e;
    FD1S1A next_ack_flag_I_0 (.D(next_addr_7__N_1160[6]), .CK(next_ack_flag_N_1498), 
           .Q(next_ack_flag)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(231[5] 1039[8])
    defparam next_ack_flag_I_0.GSR = "DISABLED";
    FD1S1D i19953 (.D(n53885), .CK(byte_rd_left_5__N_1265), .CD(byte_rd_left_5__N_1279), 
           .Q(n30625));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(225[14] 227[12])
    defparam i19953.GSR = "DISABLED";
    FD1S3DX byte_rd_left_i2 (.D(byte_rd_left_5__N_1248[2]), .CK(data_latch), 
            .CD(byte_rd_left_5__N_1255), .Q(byte_rd_left[2])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(225[14] 227[12])
    defparam byte_rd_left_i2.GSR = "DISABLED";
    LUT4 i26772_4_lut_4_lut (.A(n52425), .B(data_latch), .C(\i2c_top_debug[0] ), 
         .D(next_data_latch_N_1505), .Z(n32)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(976[30:91])
    defparam i26772_4_lut_4_lut.init = 16'hc0e0;
    LUT4 mux_464_Mux_2_i25_4_lut (.A(n52466), .B(n52241), .C(\i2c_top_debug[1] ), 
         .D(n4_adj_5203), .Z(n25)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam mux_464_Mux_2_i25_4_lut.init = 16'hc5c0;
    LUT4 n53177_bdd_3_lut_4_lut (.A(n51536), .B(\i2c_top_debug[5] ), .C(\i2c_top_debug[2] ), 
         .D(n53177), .Z(n53178)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A (C+!(D)))) */ ;
    defparam n53177_bdd_3_lut_4_lut.init = 16'h2f20;
    LUT4 n49498_bdd_3_lut_41277_then_4_lut (.A(n52425), .B(data_latch), 
         .C(n7628), .D(\i2c_top_debug[0] ), .Z(n53882)) /* synthesis lut_function=(!(A (B (C+(D))+!B (D))+!A !(((D)+!C)+!B))) */ ;
    defparam n49498_bdd_3_lut_41277_then_4_lut.init = 16'h553f;
    PFUMX i38664 (.BLUT(n21941), .ALUT(n21), .C0(n53886), .Z(n49459));
    LUT4 i26208_4_lut_4_lut (.A(n52193), .B(n63), .C(n77[5]), .D(count_wd_delay[5]), 
         .Z(count_wd_delay_31__N_1216[5])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[19:72])
    defparam i26208_4_lut_4_lut.init = 16'h5140;
    LUT4 i2c_top_debug_0__bdd_4_lut_41024 (.A(\i2c_top_debug[0] ), .B(n48117), 
         .C(n15), .D(\i2c_top_debug[4] ), .Z(n52142)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;
    defparam i2c_top_debug_0__bdd_4_lut_41024.init = 16'h77f0;
    PFUMX i2c_top_debug_5__I_0_767_Mux_1_i31 (.BLUT(n49064), .ALUT(n30_adj_5204), 
          .C0(\i2c_top_debug[4] ), .Z(n31_adj_5205)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;
    LUT4 i19952_3_lut_rep_503 (.A(n30623), .B(n30622), .C(n30621), .Z(n52439)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(225[14] 227[12])
    defparam i19952_3_lut_rep_503.init = 16'h3535;
    LUT4 i7651_2_lut_rep_350_4_lut (.A(n30623), .B(n30622), .C(n30621), 
         .D(byte_rd_left[1]), .Z(n52286)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(225[14] 227[12])
    defparam i7651_2_lut_rep_350_4_lut.init = 16'hffca;
    LUT4 i40500_then_4_lut (.A(\i2c_top_debug[0] ), .B(\i2c_top_debug[1] ), 
         .C(n32988), .D(n52425), .Z(n52607)) /* synthesis lut_function=(!(A (B (D)+!B !(C))+!A !(B))) */ ;
    defparam i40500_then_4_lut.init = 16'h64ec;
    LUT4 i40500_else_4_lut (.A(\i2c_top_debug[0] ), .B(n47361), .C(\i2c_top_debug[1] ), 
         .D(n32988), .Z(n52606)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (C)) */ ;
    defparam i40500_else_4_lut.init = 16'hdad0;
    LUT4 i2_3_lut (.A(n4068), .B(read_action), .C(write_action), .Z(n47361)) /* synthesis lut_function=((B+!(C))+!A) */ ;
    defparam i2_3_lut.init = 16'hdfdf;
    PFUMX i2c_top_debug_5__I_0_767_Mux_6_i31 (.BLUT(n15_adj_5206), .ALUT(n18960), 
          .C0(\i2c_top_debug[4] ), .Z(n31_adj_5207)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;
    LUT4 i1_2_lut_4_lut (.A(n30623), .B(n30622), .C(n30621), .D(byte_rd_left[1]), 
         .Z(byte_rd_left_5__N_1248[1])) /* synthesis lut_function=(A (B (D)+!B !(C (D)+!C !(D)))+!A (B (C (D)+!C !(D))+!B !(D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(225[14] 227[12])
    defparam i1_2_lut_4_lut.init = 16'hca35;
    LUT4 n53172_bdd_2_lut (.A(n53172), .B(\i2c_top_debug[5] ), .Z(n53173)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam n53172_bdd_2_lut.init = 16'h2222;
    LUT4 n49498_bdd_3_lut (.A(n49498), .B(n53883), .C(\i2c_top_debug[2] ), 
         .Z(n53171)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n49498_bdd_3_lut.init = 16'hcaca;
    LUT4 i26209_4_lut_4_lut (.A(n52193), .B(n63), .C(n77[4]), .D(count_wd_delay[4]), 
         .Z(count_wd_delay_31__N_1216[4])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[19:72])
    defparam i26209_4_lut_4_lut.init = 16'h5140;
    FD1S1I next_data_tx_7__I_0_i2 (.D(n51768), .CK(next_addr_7__N_1168), 
           .CD(\i2c_top_debug[5] ), .Q(next_data_tx[1])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(231[5] 1039[8])
    defparam next_data_tx_7__I_0_i2.GSR = "DISABLED";
    FD1S1I next_data_tx_7__I_0_i3 (.D(n51856), .CK(next_addr_7__N_1168), 
           .CD(\i2c_top_debug[5] ), .Q(next_data_tx[2])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(231[5] 1039[8])
    defparam next_data_tx_7__I_0_i3.GSR = "DISABLED";
    FD1S1I next_data_tx_7__I_0_i4 (.D(n51924), .CK(next_addr_7__N_1168), 
           .CD(\i2c_top_debug[5] ), .Q(next_data_tx[3])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(231[5] 1039[8])
    defparam next_data_tx_7__I_0_i4.GSR = "DISABLED";
    FD1S1I next_data_tx_7__I_0_i5 (.D(n49440), .CK(next_addr_7__N_1168), 
           .CD(\i2c_top_debug[5] ), .Q(next_data_tx[4])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(231[5] 1039[8])
    defparam next_data_tx_7__I_0_i5.GSR = "DISABLED";
    FD1S1I next_data_tx_7__I_0_i6 (.D(n51741), .CK(next_addr_7__N_1168), 
           .CD(\i2c_top_debug[5] ), .Q(next_data_tx[5])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(231[5] 1039[8])
    defparam next_data_tx_7__I_0_i6.GSR = "DISABLED";
    FD1S1I next_data_tx_7__I_0_i7 (.D(n45689), .CK(next_addr_7__N_1168), 
           .CD(\i2c_top_debug[5] ), .Q(next_data_tx[6])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(231[5] 1039[8])
    defparam next_data_tx_7__I_0_i7.GSR = "DISABLED";
    FD1S1I next_data_tx_7__I_0_i8 (.D(n49392), .CK(next_addr_7__N_1168), 
           .CD(\i2c_top_debug[5] ), .Q(next_data_tx[7])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(231[5] 1039[8])
    defparam next_data_tx_7__I_0_i8.GSR = "DISABLED";
    FD1S1A next_addr_7__I_0_i2 (.D(next_addr_7__N_1160[1]), .CK(next_addr_7__N_1168), 
           .Q(next_addr[1])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(231[5] 1039[8])
    defparam next_addr_7__I_0_i2.GSR = "DISABLED";
    FD1S1A next_addr_7__I_0_i3 (.D(next_addr_7__N_1160[2]), .CK(next_addr_7__N_1168), 
           .Q(next_addr[2])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(231[5] 1039[8])
    defparam next_addr_7__I_0_i3.GSR = "DISABLED";
    LUT4 data_latch_I_0_772_2_lut (.A(data_latch), .B(one_byte_ready), .Z(module_data_out_7__N_1332)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(209[18:66])
    defparam data_latch_I_0_772_2_lut.init = 16'h2222;
    LUT4 i26194_4_lut_4_lut (.A(n52193), .B(n63), .C(n77[8]), .D(count_wd_delay[8]), 
         .Z(count_wd_delay_31__N_1216[8])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[19:72])
    defparam i26194_4_lut_4_lut.init = 16'h5140;
    LUT4 i4_4_lut (.A(n52452), .B(\i2c_top_debug[4] ), .C(\i2c_top_debug[1] ), 
         .D(\i2c_top_debug[5] ), .Z(resetn_imu_N_1182)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i4_4_lut.init = 16'hfffe;
    PFUMX i38607 (.BLUT(n10_adj_5208), .ALUT(n6), .C0(\next_i2c_device_driver_state[3] ), 
          .Z(n49402));
    PFUMX i38608 (.BLUT(n46519), .ALUT(n46521), .C0(\next_i2c_device_driver_state[3] ), 
          .Z(n49403));
    LUT4 i26168_4_lut_4_lut (.A(n52193), .B(n63), .C(n77[30]), .D(count_wd_delay[30]), 
         .Z(count_wd_delay_31__N_1216[30])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[19:72])
    defparam i26168_4_lut_4_lut.init = 16'h5140;
    LUT4 n51918_bdd_4_lut (.A(n51918), .B(n51917), .C(\i2c_top_debug[3] ), 
         .D(\i2c_top_debug[2] ), .Z(n53875)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam n51918_bdd_4_lut.init = 16'hca00;
    LUT4 i2c_top_debug_0__bdd_4_lut_40715 (.A(\i2c_top_debug[0] ), .B(\i2c_top_debug[1] ), 
         .C(\data_reg[5] ), .D(n52228), .Z(n51738)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2c_top_debug_0__bdd_4_lut_40715.init = 16'h8000;
    LUT4 n51740_bdd_3_lut (.A(n51740), .B(n53872), .C(\i2c_top_debug[4] ), 
         .Z(n51741)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n51740_bdd_3_lut.init = 16'hcaca;
    LUT4 i33211_4_lut_4_lut_4_lut (.A(data_rx_adj_5257[6]), .B(\i2c_top_debug[3] ), 
         .C(n4_adj_5210), .D(n52425), .Z(n43987)) /* synthesis lut_function=(A (B (C)+!B !(D))+!A (B+!(D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1010[28:70])
    defparam i33211_4_lut_4_lut_4_lut.init = 16'hc4f7;
    LUT4 i1_2_lut_4_lut_adj_282 (.A(n52205), .B(n52289), .C(n52288), .D(n63), 
         .Z(sys_clk_enable_231)) /* synthesis lut_function=((B (D)+!B ((D)+!C))+!A) */ ;
    defparam i1_2_lut_4_lut_adj_282.init = 16'hff57;
    LUT4 i1_2_lut_rep_252_3_lut_4_lut (.A(\i2c_top_debug[1] ), .B(n52306), 
         .C(n66), .D(n52318), .Z(n52188)) /* synthesis lut_function=(A (C+(D))+!A ((C+(D))+!B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i1_2_lut_rep_252_3_lut_4_lut.init = 16'hfff1;
    FD1S3IX wd_event_active_687 (.D(n52174), .CK(sys_clk), .CD(n63), .Q(wd_event_active)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[14] 151[12])
    defparam wd_event_active_687.GSR = "ENABLED";
    FD1S3IX data_latch_694 (.D(n2486[5]), .CK(sys_clk), .CD(wd_event_active), 
            .Q(data_latch)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam data_latch_694.GSR = "ENABLED";
    LUT4 n28056_bdd_4_lut_40656 (.A(n52200), .B(\i2c_top_debug[3] ), .C(\data_reg[1] ), 
         .D(\i2c_top_debug[1] ), .Z(n51764)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam n28056_bdd_4_lut_40656.init = 16'h2000;
    LUT4 n10_bdd_4_lut (.A(n10), .B(n14), .C(\i2c_top_debug[2] ), .D(\i2c_top_debug[3] ), 
         .Z(n51767)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C+!(D)))) */ ;
    defparam n10_bdd_4_lut.init = 16'hcacc;
    LUT4 n51767_bdd_3_lut (.A(n51767), .B(n51766), .C(\i2c_top_debug[4] ), 
         .Z(n51768)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n51767_bdd_3_lut.init = 16'hcaca;
    LUT4 i7659_2_lut_rep_303_3_lut (.A(byte_rd_left[1]), .B(n52439), .C(byte_rd_left[2]), 
         .Z(n52239)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(226[29:50])
    defparam i7659_2_lut_rep_303_3_lut.init = 16'hfbfb;
    LUT4 i1_2_lut (.A(data_rx_adj_5257[2]), .B(data_rx_adj_5257[4]), .Z(n1516)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut.init = 16'h4444;
    LUT4 i39162_1_lut_3_lut (.A(n19779), .B(n38357), .C(\i2c_top_debug[5] ), 
         .Z(n49768)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i39162_1_lut_3_lut.init = 16'h3535;
    LUT4 i1_2_lut_3_lut (.A(byte_rd_left[1]), .B(n52439), .C(byte_rd_left[2]), 
         .Z(byte_rd_left_5__N_1248[2])) /* synthesis lut_function=(A (C)+!A !(B (C)+!B !(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(226[29:50])
    defparam i1_2_lut_3_lut.init = 16'hb4b4;
    LUT4 i1_2_lut_3_lut_4_lut_rep_351 (.A(byte_rd_left[1]), .B(n52439), 
         .C(byte_rd_left[3]), .D(byte_rd_left[2]), .Z(n52287)) /* synthesis lut_function=(A (C)+!A (B (C (D)+!C !(D))+!B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(226[29:50])
    defparam i1_2_lut_3_lut_4_lut_rep_351.init = 16'hf0b4;
    LUT4 i4_4_lut_4_lut (.A(byte_rd_left[1]), .B(n52439), .C(byte_rd_left[3]), 
         .D(byte_rd_left[2]), .Z(n10_adj_5212)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(226[29:50])
    defparam i4_4_lut_4_lut.init = 16'h0001;
    LUT4 i1_3_lut_4_lut (.A(\i2c_top_debug[5] ), .B(n52464), .C(next_addr_7__N_1168), 
         .D(n26115), .Z(next_ack_flag_N_1498)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i1_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i2c_top_debug_1__bdd_4_lut_40633 (.A(\i2c_top_debug[1] ), .B(\i2c_top_debug[0] ), 
         .C(n52425), .D(data_rx_adj_5257[6]), .Z(n50986)) /* synthesis lut_function=(A (B (C)+!B !((D)+!C))) */ ;
    defparam i2c_top_debug_1__bdd_4_lut_40633.init = 16'h80a0;
    LUT4 i26212_4_lut_4_lut (.A(n52193), .B(n63), .C(n77[3]), .D(count_wd_delay[3]), 
         .Z(count_wd_delay_31__N_1216[3])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[19:72])
    defparam i26212_4_lut_4_lut.init = 16'h5140;
    LUT4 i33673_2_lut (.A(byte_wr_left[1]), .B(byte_wr_left[0]), .Z(n2[1])) /* synthesis lut_function=(A (B)+!A !(B)) */ ;
    defparam i33673_2_lut.init = 16'h9999;
    LUT4 i1_2_lut_adj_283 (.A(is_2_byte_reg), .B(n48107), .Z(n48108)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[14] 151[12])
    defparam i1_2_lut_adj_283.init = 16'h8888;
    LUT4 i27604_3_lut_4_lut (.A(\i2c_top_debug[2] ), .B(n52425), .C(\i2c_top_debug[1] ), 
         .D(\i2c_top_debug[0] ), .Z(n29_adj_5214)) /* synthesis lut_function=(!(A+(B+(C (D)+!C !(D))))) */ ;
    defparam i27604_3_lut_4_lut.init = 16'h0110;
    PFUMX i15786 (.BLUT(n26203), .ALUT(n26271), .C0(\i2c_top_debug[3] ), 
          .Z(n26272));
    LUT4 byte_rd_left_5__N_1255_I_0_757_2_lut (.A(byte_rd_left_5__N_1255), 
         .B(\target_read_count[0] ), .Z(byte_rd_left_5__N_1266)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(225[14] 227[12])
    defparam byte_rd_left_5__N_1255_I_0_757_2_lut.init = 16'h8888;
    LUT4 i39642_2_lut (.A(byte_rd_left_5__N_1255), .B(\target_read_count[0] ), 
         .Z(byte_rd_left_5__N_1282)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i39642_2_lut.init = 16'h2222;
    LUT4 i2c_top_debug_0__bdd_4_lut_40758 (.A(\i2c_top_debug[0] ), .B(\i2c_top_debug[1] ), 
         .C(\data_reg[2] ), .D(n52228), .Z(n51853)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2c_top_debug_0__bdd_4_lut_40758.init = 16'h8000;
    LUT4 i27562_4_lut (.A(n4068), .B(n52424), .C(write_action), .D(read_action), 
         .Z(n6_c)) /* synthesis lut_function=(!(A (B (C+(D))))) */ ;
    defparam i27562_4_lut.init = 16'h777f;
    LUT4 i38593_4_lut (.A(n52263), .B(n50), .C(\i2c_top_debug[2] ), .D(n52293), 
         .Z(n49388)) /* synthesis lut_function=(!(A (B (C (D)))+!A (B ((D)+!C)+!B !(C)))) */ ;
    defparam i38593_4_lut.init = 16'h3afa;
    LUT4 i1_2_lut_adj_284 (.A(\i2c_top_debug[2] ), .B(\i2c_top_debug[0] ), 
         .Z(n48025)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i1_2_lut_adj_284.init = 16'h2222;
    LUT4 i25795_4_lut (.A(count_wd_delay[0]), .B(n52193), .C(n77[0]), 
         .D(n63), .Z(count_wd_delay_31__N_1216[0])) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(144[14] 151[12])
    defparam i25795_4_lut.init = 16'h3022;
    LUT4 i39894_4_lut (.A(n49), .B(n62), .C(n58), .D(n50_adj_5215), 
         .Z(n63)) /* synthesis lut_function=(!(A (B (C (D))))) */ ;
    defparam i39894_4_lut.init = 16'h7fff;
    LUT4 i17_4_lut (.A(count_wd_delay[0]), .B(count_wd_delay[10]), .C(count_wd_delay[27]), 
         .D(count_wd_delay[25]), .Z(n49)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i17_4_lut.init = 16'h8000;
    LUT4 i30_4_lut (.A(n41), .B(n60), .C(n54), .D(n42), .Z(n62)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i30_4_lut.init = 16'h8000;
    LUT4 i26_4_lut (.A(count_wd_delay[3]), .B(n52), .C(n38), .D(count_wd_delay[15]), 
         .Z(n58)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i26_4_lut.init = 16'h8000;
    LUT4 i18_4_lut (.A(count_wd_delay[29]), .B(count_wd_delay[17]), .C(count_wd_delay[19]), 
         .D(count_wd_delay[8]), .Z(n50_adj_5215)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i18_4_lut.init = 16'h8000;
    LUT4 i9_2_lut (.A(count_wd_delay[31]), .B(count_wd_delay[13]), .Z(n41)) /* synthesis lut_function=(A (B)) */ ;
    defparam i9_2_lut.init = 16'h8888;
    FD1S3IX i2c_cmd_state__i6 (.D(next_i2c_cmd_state_5__N_1479[5]), .CK(sys_clk), 
            .CD(wd_event_active), .Q(\i2c_top_debug[5] )) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam i2c_cmd_state__i6.GSR = "ENABLED";
    LUT4 i28_4_lut (.A(count_wd_delay[4]), .B(n56), .C(n46), .D(count_wd_delay[24]), 
         .Z(n60)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i28_4_lut.init = 16'h8000;
    LUT4 n1304_bdd_4_lut_40897 (.A(n1296[0]), .B(\i2c_top_debug[2] ), .C(data_tx[0]), 
         .D(\i2c_top_debug[0] ), .Z(n51003)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A (((D)+!C)+!B))) */ ;
    defparam n1304_bdd_4_lut_40897.init = 16'h22c0;
    LUT4 i22_4_lut (.A(count_wd_delay[6]), .B(count_wd_delay[14]), .C(count_wd_delay[22]), 
         .D(count_wd_delay[30]), .Z(n54)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i22_4_lut.init = 16'h8000;
    PFUMX mux_464_Mux_0_i25 (.BLUT(n37968), .ALUT(n24_adj_5217), .C0(\i2c_top_debug[1] ), 
          .Z(n25_adj_5218)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;
    LUT4 i10_2_lut (.A(count_wd_delay[23]), .B(count_wd_delay[20]), .Z(n42)) /* synthesis lut_function=(A (B)) */ ;
    defparam i10_2_lut.init = 16'h8888;
    LUT4 i24_4_lut (.A(count_wd_delay[21]), .B(count_wd_delay[2]), .C(count_wd_delay[16]), 
         .D(count_wd_delay[28]), .Z(n56)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i24_4_lut.init = 16'h8000;
    LUT4 i14_2_lut (.A(count_wd_delay[12]), .B(count_wd_delay[26]), .Z(n46)) /* synthesis lut_function=(A (B)) */ ;
    defparam i14_2_lut.init = 16'h8888;
    LUT4 i20_4_lut (.A(count_wd_delay[1]), .B(count_wd_delay[11]), .C(count_wd_delay[9]), 
         .D(count_wd_delay[18]), .Z(n52)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i20_4_lut.init = 16'h8000;
    FD1S3IX i2c_cmd_state__i5 (.D(n49419), .CK(sys_clk), .CD(n37653), 
            .Q(\i2c_top_debug[4] )) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam i2c_cmd_state__i5.GSR = "ENABLED";
    FD1S3IX i2c_cmd_state__i4 (.D(n49395), .CK(sys_clk), .CD(n37653), 
            .Q(\i2c_top_debug[3] )) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam i2c_cmd_state__i4.GSR = "ENABLED";
    FD1S3IX i2c_cmd_state__i3 (.D(next_i2c_cmd_state_5__N_1479[2]), .CK(sys_clk), 
            .CD(wd_event_active), .Q(\i2c_top_debug[2] )) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam i2c_cmd_state__i3.GSR = "ENABLED";
    FD1S3IX i2c_cmd_state__i2 (.D(next_i2c_cmd_state_5__N_1479[1]), .CK(sys_clk), 
            .CD(wd_event_active), .Q(\i2c_top_debug[1] )) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam i2c_cmd_state__i2.GSR = "ENABLED";
    LUT4 mux_464_Mux_0_i21_4_lut_4_lut (.A(data_rx_adj_5257[2]), .B(n52425), 
         .C(\i2c_top_debug[0] ), .D(\i2c_top_debug[1] ), .Z(n21)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B (C (D))+!B !(C)))) */ ;
    defparam mux_464_Mux_0_i21_4_lut_4_lut.init = 16'h3c7c;
    LUT4 i6_2_lut (.A(count_wd_delay[5]), .B(count_wd_delay[7]), .Z(n38)) /* synthesis lut_function=(A (B)) */ ;
    defparam i6_2_lut.init = 16'h8888;
    LUT4 i2_3_lut_4_lut (.A(data_rx_adj_5257[2]), .B(n52425), .C(n37653), 
         .D(n27391), .Z(n48107)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;
    defparam i2_3_lut_4_lut.init = 16'h0800;
    LUT4 i2c_top_debug_0__bdd_4_lut_40899 (.A(\i2c_top_debug[0] ), .B(\i2c_top_debug[1] ), 
         .C(\data_reg[3] ), .D(n52228), .Z(n51921)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2c_top_debug_0__bdd_4_lut_40899.init = 16'h8000;
    LUT4 i25450_4_lut_4_lut (.A(n52425), .B(\data_reg[4] ), .C(\i2c_top_debug[1] ), 
         .D(n27301), .Z(n10_adj_5219)) /* synthesis lut_function=(A (B (C (D)))+!A (B ((D)+!C)+!B !(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i25450_4_lut_4_lut.init = 16'hc505;
    LUT4 read_write_in_I_0_1_lut (.A(read_write_in), .Z(read_write_in_N_1023)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(830[24:50])
    defparam read_write_in_I_0_1_lut.init = 16'h5555;
    LUT4 i1_4_lut_4_lut (.A(n52425), .B(\i2c_top_debug[0] ), .C(\i2c_top_debug[1] ), 
         .D(n12), .Z(n46343)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i1_4_lut_4_lut.init = 16'h5140;
    LUT4 i19956_3_lut (.A(n30627), .B(n30626), .C(n30625), .Z(byte_rd_left[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(225[14] 227[12])
    defparam i19956_3_lut.init = 16'hcaca;
    LUT4 i2c_top_debug_5__I_0_767_Mux_2_i28_4_lut_4_lut_4_lut (.A(n52425), 
         .B(data_latch), .C(\i2c_top_debug[1] ), .D(\i2c_top_debug[0] ), 
         .Z(n28)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A (B (C+!(D))+!B (C (D)+!C !(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i2c_top_debug_5__I_0_767_Mux_2_i28_4_lut_4_lut_4_lut.init = 16'h0530;
    LUT4 i2c_top_debug_5__I_0_767_Mux_6_i63_3_lut (.A(n31_adj_5207), .B(n38357), 
         .C(\i2c_top_debug[5] ), .Z(next_addr_7__N_1160[6])) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i2c_top_debug_5__I_0_767_Mux_6_i63_3_lut.init = 16'h3a3a;
    LUT4 i27637_4_lut (.A(n52425), .B(n27058), .C(n48426), .D(\i2c_top_debug[0] ), 
         .Z(n38357)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A ((C (D))+!B)) */ ;
    defparam i27637_4_lut.init = 16'hf3bb;
    LUT4 i37640_2_lut (.A(\i2c_top_debug[1] ), .B(data_latch), .Z(n48426)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i37640_2_lut.init = 16'heeee;
    LUT4 n7_bdd_3_lut_40761_4_lut_4_lut (.A(n52425), .B(n51854), .C(\i2c_top_debug[3] ), 
         .D(n52273), .Z(n51855)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam n7_bdd_3_lut_40761_4_lut_4_lut.init = 16'hc5c0;
    LUT4 i1_4_lut_4_lut_adj_285 (.A(n52425), .B(\i2c_top_debug[0] ), .C(\i2c_top_debug[1] ), 
         .D(\i2c_top_debug[2] ), .Z(n49_adj_5220)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i1_4_lut_4_lut_adj_285.init = 16'h5140;
    LUT4 n7_bdd_3_lut_40653_4_lut_4_lut (.A(n52425), .B(n51739), .C(\i2c_top_debug[3] ), 
         .D(n52273), .Z(n51740)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam n7_bdd_3_lut_40653_4_lut_4_lut.init = 16'hc5c0;
    LUT4 byte_rd_left_5__N_1255_I_0_756_2_lut (.A(byte_rd_left_5__N_1255), 
         .B(\target_read_count[1] ), .Z(byte_rd_left_5__N_1265)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(225[14] 227[12])
    defparam byte_rd_left_5__N_1255_I_0_756_2_lut.init = 16'h8888;
    LUT4 i2_3_lut_3_lut_4_lut (.A(\i2c_top_debug[3] ), .B(\i2c_top_debug[0] ), 
         .C(\i2c_top_debug[1] ), .D(\i2c_top_debug[2] ), .Z(n48722)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(267[14] 1038[12])
    defparam i2_3_lut_3_lut_4_lut.init = 16'h0020;
    LUT4 i39640_2_lut (.A(byte_rd_left_5__N_1255), .B(\target_read_count[1] ), 
         .Z(byte_rd_left_5__N_1279)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i39640_2_lut.init = 16'h2222;
    LUT4 i26213_4_lut_4_lut (.A(n52193), .B(n63), .C(n77[2]), .D(count_wd_delay[2]), 
         .Z(count_wd_delay_31__N_1216[2])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[19:72])
    defparam i26213_4_lut_4_lut.init = 16'h5140;
    LUT4 n7_bdd_3_lut_4_lut_4_lut (.A(n52425), .B(n51922), .C(\i2c_top_debug[3] ), 
         .D(n52273), .Z(n51923)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam n7_bdd_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 i37609_4_lut_4_lut (.A(n52425), .B(\i2c_top_debug[4] ), .C(n52424), 
         .D(n9), .Z(n48394)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i37609_4_lut_4_lut.init = 16'h5140;
    LUT4 i15723_2_lut_3_lut_3_lut (.A(\i2c_top_debug[1] ), .B(\i2c_top_debug[2] ), 
         .C(\i2c_top_debug[0] ), .Z(n26203)) /* synthesis lut_function=(!(A (B (C)+!B !(C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam i15723_2_lut_3_lut_3_lut.init = 16'h7d7d;
    LUT4 i27290_4_lut_4_lut (.A(n52425), .B(n52466), .C(\i2c_top_debug[0] ), 
         .D(n52459), .Z(n37968)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A !(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i27290_4_lut_4_lut.init = 16'h5052;
    LUT4 mux_464_Mux_1_i23_4_lut_4_lut (.A(n52425), .B(n52466), .C(\i2c_top_debug[0] ), 
         .D(n52459), .Z(n23)) /* synthesis lut_function=(A (B (C)+!B (C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam mux_464_Mux_1_i23_4_lut_4_lut.init = 16'ha2a0;
    LUT4 i38724_4_lut (.A(\i2c_top_debug[1] ), .B(n32988), .C(\i2c_top_debug[0] ), 
         .D(n5), .Z(n49519)) /* synthesis lut_function=(!(A (C (D))+!A !(B (C)))) */ ;
    defparam i38724_4_lut.init = 16'h4aea;
    LUT4 n15_bdd_3_lut (.A(n28), .B(n38357), .C(\i2c_top_debug[5] ), .Z(n52024)) /* synthesis lut_function=(!(A (B (C))+!A (B+!(C)))) */ ;
    defparam n15_bdd_3_lut.init = 16'h3a3a;
    LUT4 i26956_4_lut_4_lut_4_lut (.A(\i2c_top_debug[1] ), .B(n48), .C(n27058), 
         .D(\i2c_top_debug[0] ), .Z(n62_adj_5221)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A !(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam i26956_4_lut_4_lut_4_lut.init = 16'h50d0;
    LUT4 i26054_rep_312_4_lut (.A(\i2c_top_debug[5] ), .B(n52464), .C(n53886), 
         .D(\i2c_top_debug[1] ), .Z(n52248)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i26054_rep_312_4_lut.init = 16'hfffe;
    LUT4 i26214_4_lut_4_lut (.A(n52193), .B(n63), .C(n77[1]), .D(count_wd_delay[1]), 
         .Z(count_wd_delay_31__N_1216[1])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[19:72])
    defparam i26214_4_lut_4_lut.init = 16'h5140;
    LUT4 i1_4_lut (.A(\i2c_top_debug[1] ), .B(n52234), .C(n33015), .D(\i2c_top_debug[0] ), 
         .Z(n22)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (B+(C (D)))) */ ;
    defparam i1_4_lut.init = 16'hfcee;
    LUT4 i1_4_lut_4_lut_adj_286 (.A(\i2c_top_debug[1] ), .B(\data_reg[4] ), 
         .C(n52455), .D(n53886), .Z(n12)) /* synthesis lut_function=(A (B (C (D)))+!A (D)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam i1_4_lut_4_lut_adj_286.init = 16'hd500;
    LUT4 i38666_3_lut (.A(n49459), .B(n49460), .C(\i2c_top_debug[3] ), 
         .Z(n49461)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38666_3_lut.init = 16'hcaca;
    LUT4 i14085_2_lut_rep_380 (.A(\i2c_top_debug[0] ), .B(\i2c_top_debug[1] ), 
         .Z(n52316)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i14085_2_lut_rep_380.init = 16'hbbbb;
    LUT4 i1_2_lut_3_lut_adj_287 (.A(\i2c_top_debug[0] ), .B(\i2c_top_debug[1] ), 
         .C(data_tx[6]), .Z(n9)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i1_2_lut_3_lut_adj_287.init = 16'h4040;
    LUT4 i27086_2_lut_3_lut_4_lut (.A(\i2c_top_debug[0] ), .B(\i2c_top_debug[1] ), 
         .C(n52425), .D(\i2c_top_debug[2] ), .Z(n29_adj_5202)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i27086_2_lut_3_lut_4_lut.init = 16'h0004;
    LUT4 i1_2_lut_3_lut_4_lut (.A(\i2c_top_debug[0] ), .B(\i2c_top_debug[1] ), 
         .C(n1296[0]), .D(n52425), .Z(n4)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0040;
    LUT4 i2c_top_debug_0__bdd_2_lut_3_lut_4_lut (.A(\i2c_top_debug[0] ), .B(\i2c_top_debug[1] ), 
         .C(data_tx[2]), .D(n52425), .Z(n51852)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i2c_top_debug_0__bdd_2_lut_3_lut_4_lut.init = 16'h0040;
    LUT4 n27301_bdd_2_lut_3_lut_4_lut (.A(\i2c_top_debug[0] ), .B(\i2c_top_debug[1] ), 
         .C(data_tx[3]), .D(n52425), .Z(n51759)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam n27301_bdd_2_lut_3_lut_4_lut.init = 16'h0040;
    LUT4 i2c_top_debug_0__bdd_2_lut_40714_3_lut_4_lut (.A(\i2c_top_debug[0] ), 
         .B(\i2c_top_debug[1] ), .C(data_tx[5]), .D(n52425), .Z(n51737)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i2c_top_debug_0__bdd_2_lut_40714_3_lut_4_lut.init = 16'h0040;
    LUT4 i12563_3_lut_4_lut (.A(\i2c_top_debug[0] ), .B(\i2c_top_debug[1] ), 
         .C(n52425), .D(data_latch), .Z(n19779)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i12563_3_lut_4_lut.init = 16'hf4b0;
    LUT4 i38723_4_lut_4_lut (.A(\i2c_top_debug[1] ), .B(n4_adj_5222), .C(\i2c_top_debug[5] ), 
         .D(n49516), .Z(n49518)) /* synthesis lut_function=(!(A (C+!(D))+!A !(B (C+(D))+!B !(C+!(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam i38723_4_lut_4_lut.init = 16'h4f40;
    FD1S3AX data_tx_i7 (.D(next_data_tx[7]), .CK(sys_clk), .Q(data_tx_c[7])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam data_tx_i7.GSR = "ENABLED";
    FD1S3AX data_tx_i6 (.D(next_data_tx[6]), .CK(sys_clk), .Q(data_tx_c[6])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam data_tx_i6.GSR = "ENABLED";
    FD1S3AX data_tx_i5 (.D(next_data_tx[5]), .CK(sys_clk), .Q(data_tx_c[5])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam data_tx_i5.GSR = "ENABLED";
    FD1S3AX data_tx_i4 (.D(next_data_tx[4]), .CK(sys_clk), .Q(data_tx_c[4])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam data_tx_i4.GSR = "ENABLED";
    FD1S3AX data_tx_i3 (.D(next_data_tx[3]), .CK(sys_clk), .Q(data_tx_c[3])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam data_tx_i3.GSR = "ENABLED";
    FD1S3AX data_tx_i2 (.D(next_data_tx[2]), .CK(sys_clk), .Q(data_tx_c[2])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam data_tx_i2.GSR = "ENABLED";
    FD1S3AX data_tx_i1 (.D(next_data_tx[1]), .CK(sys_clk), .Q(data_tx_c[1])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam data_tx_i1.GSR = "ENABLED";
    FD1S3AX addr_i3 (.D(next_addr[2]), .CK(sys_clk), .Q(addr[2])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam addr_i3.GSR = "ENABLED";
    FD1S3AX addr_i2 (.D(next_addr[1]), .CK(sys_clk), .Q(addr[1])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam addr_i2.GSR = "ENABLED";
    LUT4 i10_4_lut_4_lut (.A(\i2c_top_debug[1] ), .B(\i2c_top_debug[3] ), 
         .C(n52425), .D(count_us_11__N_1299), .Z(n8)) /* synthesis lut_function=(!(A (B (C)+!B (D))+!A (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam i10_4_lut_4_lut.init = 16'h0d2f;
    FD1S3AY count_us_i0_i10_19926_19927_set (.D(n26[10]), .CK(sys_clk), 
            .Q(n30598)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(128[14] 131[34])
    defparam count_us_i0_i10_19926_19927_set.GSR = "ENABLED";
    LUT4 i1_4_lut_adj_288 (.A(n27058), .B(n52299), .C(n12368[0]), .D(\i2c_top_debug[0] ), 
         .Z(n4_adj_5222)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))) */ ;
    defparam i1_4_lut_adj_288.init = 16'ha022;
    LUT4 i5_4_lut (.A(n52286), .B(byte_rd_left[3]), .C(n8_adj_5228), .D(byte_rd_left[2]), 
         .Z(next_data_latch_N_1505)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(982[28:49])
    defparam i5_4_lut.init = 16'hfffe;
    FD1S3AY count_us_i0_i9_19929_19930_set (.D(n26[9]), .CK(sys_clk), .Q(n30601)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(128[14] 131[34])
    defparam count_us_i0_i9_19929_19930_set.GSR = "ENABLED";
    FD1S3AY count_us_i0_i8_19932_19933_set (.D(n26[8]), .CK(sys_clk), .Q(n30604)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(128[14] 131[34])
    defparam count_us_i0_i8_19932_19933_set.GSR = "ENABLED";
    LUT4 i2_2_lut (.A(byte_rd_left[5]), .B(byte_rd_left[4]), .Z(n8_adj_5228)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(982[28:49])
    defparam i2_2_lut.init = 16'heeee;
    FD1S3AY count_us_i0_i6_19935_19936_set (.D(n26[6]), .CK(sys_clk), .Q(n30607)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(128[14] 131[34])
    defparam count_us_i0_i6_19935_19936_set.GSR = "ENABLED";
    FD1P3BX count_us_i0_i7 (.D(count_us_11__N_1287[7]), .SP(count_us_11__N_1299), 
            .CK(sys_clk), .PD(count_us_11__N_1209), .Q(count_us[7])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(128[14] 131[34])
    defparam count_us_i0_i7.GSR = "DISABLED";
    FD1S3AY count_us_i0_i0_19938_19939_set (.D(n26[0]), .CK(sys_clk), .Q(n30610)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(128[14] 131[34])
    defparam count_us_i0_i0_19938_19939_set.GSR = "ENABLED";
    FD1P3BX count_us_i0_i5 (.D(count_us_11__N_1287[5]), .SP(count_us_11__N_1299), 
            .CK(sys_clk), .PD(count_us_11__N_1209), .Q(count_us[5])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(128[14] 131[34])
    defparam count_us_i0_i5.GSR = "DISABLED";
    FD1P3BX count_us_i0_i4 (.D(count_us_11__N_1287[4]), .SP(count_us_11__N_1299), 
            .CK(sys_clk), .PD(count_us_11__N_1209), .Q(count_us[4])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(128[14] 131[34])
    defparam count_us_i0_i4.GSR = "DISABLED";
    FD1P3BX count_us_i0_i3 (.D(count_us_11__N_1287[3]), .SP(count_us_11__N_1299), 
            .CK(sys_clk), .PD(count_us_11__N_1209), .Q(count_us[3])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(128[14] 131[34])
    defparam count_us_i0_i3.GSR = "DISABLED";
    LUT4 i39838_2_lut (.A(\i2c_top_debug[5] ), .B(\i2c_top_debug[4] ), .Z(n49529)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i39838_2_lut.init = 16'hbbbb;
    FD1P3BX count_us_i0_i2 (.D(count_us_11__N_1287[2]), .SP(count_us_11__N_1299), 
            .CK(sys_clk), .PD(count_us_11__N_1209), .Q(count_us[2])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(128[14] 131[34])
    defparam count_us_i0_i2.GSR = "DISABLED";
    FD1P3BX count_us_i0_i1 (.D(count_us_11__N_1287[1]), .SP(count_us_11__N_1299), 
            .CK(sys_clk), .PD(count_us_11__N_1209), .Q(count_us[1])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(128[14] 131[34])
    defparam count_us_i0_i1.GSR = "DISABLED";
    FD1P3AX module_data_out_i0_i7 (.D(data_rx_adj_5257[7]), .SP(module_data_out_7__N_1332), 
            .CK(sys_clk), .Q(data_rx[7])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(209[14] 216[12])
    defparam module_data_out_i0_i7.GSR = "ENABLED";
    FD1P3AX module_data_out_i0_i6 (.D(data_rx_adj_5257[6]), .SP(module_data_out_7__N_1332), 
            .CK(sys_clk), .Q(data_rx[6])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(209[14] 216[12])
    defparam module_data_out_i0_i6.GSR = "ENABLED";
    FD1P3AX module_data_out_i0_i5 (.D(data_rx_adj_5257[5]), .SP(module_data_out_7__N_1332), 
            .CK(sys_clk), .Q(data_rx[5])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(209[14] 216[12])
    defparam module_data_out_i0_i5.GSR = "ENABLED";
    FD1P3AX module_data_out_i0_i4 (.D(data_rx_adj_5257[4]), .SP(module_data_out_7__N_1332), 
            .CK(sys_clk), .Q(data_rx[4])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(209[14] 216[12])
    defparam module_data_out_i0_i4.GSR = "ENABLED";
    FD1P3AX module_data_out_i0_i3 (.D(data_rx_adj_5257[3]), .SP(module_data_out_7__N_1332), 
            .CK(sys_clk), .Q(data_rx[3])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(209[14] 216[12])
    defparam module_data_out_i0_i3.GSR = "ENABLED";
    FD1S3AY count_wd_delay_i31 (.D(count_wd_delay_31__N_1216[31]), .CK(sys_clk), 
            .Q(count_wd_delay[31])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[14] 151[12])
    defparam count_wd_delay_i31.GSR = "ENABLED";
    FD1P3AX module_data_out_i0_i2 (.D(data_rx_adj_5257[2]), .SP(module_data_out_7__N_1332), 
            .CK(sys_clk), .Q(data_rx[2])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(209[14] 216[12])
    defparam module_data_out_i0_i2.GSR = "ENABLED";
    FD1P3AX module_data_out_i0_i1 (.D(data_rx_adj_5257[1]), .SP(module_data_out_7__N_1332), 
            .CK(sys_clk), .Q(data_rx[1])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(209[14] 216[12])
    defparam module_data_out_i0_i1.GSR = "ENABLED";
    FD1S3AY count_wd_delay_i30 (.D(count_wd_delay_31__N_1216[30]), .CK(sys_clk), 
            .Q(count_wd_delay[30])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[14] 151[12])
    defparam count_wd_delay_i30.GSR = "ENABLED";
    FD1S3AY count_wd_delay_i29 (.D(count_wd_delay_31__N_1216[29]), .CK(sys_clk), 
            .Q(count_wd_delay[29])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[14] 151[12])
    defparam count_wd_delay_i29.GSR = "ENABLED";
    FD1S3AY count_wd_delay_i28 (.D(count_wd_delay_31__N_1216[28]), .CK(sys_clk), 
            .Q(count_wd_delay[28])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[14] 151[12])
    defparam count_wd_delay_i28.GSR = "ENABLED";
    FD1S3AY count_wd_delay_i27 (.D(count_wd_delay_31__N_1216[27]), .CK(sys_clk), 
            .Q(count_wd_delay[27])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[14] 151[12])
    defparam count_wd_delay_i27.GSR = "ENABLED";
    FD1S3AY count_wd_delay_i26 (.D(count_wd_delay_31__N_1216[26]), .CK(sys_clk), 
            .Q(count_wd_delay[26])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[14] 151[12])
    defparam count_wd_delay_i26.GSR = "ENABLED";
    FD1S3AY count_wd_delay_i25 (.D(count_wd_delay_31__N_1216[25]), .CK(sys_clk), 
            .Q(count_wd_delay[25])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[14] 151[12])
    defparam count_wd_delay_i25.GSR = "ENABLED";
    FD1S3AY count_wd_delay_i24 (.D(count_wd_delay_31__N_1216[24]), .CK(sys_clk), 
            .Q(count_wd_delay[24])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[14] 151[12])
    defparam count_wd_delay_i24.GSR = "ENABLED";
    FD1S3AY count_wd_delay_i23 (.D(count_wd_delay_31__N_1216[23]), .CK(sys_clk), 
            .Q(count_wd_delay[23])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[14] 151[12])
    defparam count_wd_delay_i23.GSR = "ENABLED";
    FD1S3AY count_wd_delay_i22 (.D(count_wd_delay_31__N_1216[22]), .CK(sys_clk), 
            .Q(count_wd_delay[22])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[14] 151[12])
    defparam count_wd_delay_i22.GSR = "ENABLED";
    FD1S3AY count_wd_delay_i20 (.D(count_wd_delay_31__N_1216[20]), .CK(sys_clk), 
            .Q(count_wd_delay[20])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[14] 151[12])
    defparam count_wd_delay_i20.GSR = "ENABLED";
    FD1S3AY count_wd_delay_i19 (.D(count_wd_delay_31__N_1216[19]), .CK(sys_clk), 
            .Q(count_wd_delay[19])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[14] 151[12])
    defparam count_wd_delay_i19.GSR = "ENABLED";
    FD1S3AY count_wd_delay_i18 (.D(count_wd_delay_31__N_1216[18]), .CK(sys_clk), 
            .Q(count_wd_delay[18])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[14] 151[12])
    defparam count_wd_delay_i18.GSR = "ENABLED";
    FD1S3AY count_wd_delay_i16 (.D(count_wd_delay_31__N_1216[16]), .CK(sys_clk), 
            .Q(count_wd_delay[16])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[14] 151[12])
    defparam count_wd_delay_i16.GSR = "ENABLED";
    LUT4 i2_2_lut_2_lut (.A(\i2c_top_debug[1] ), .B(data_rx_adj_5257[6]), 
         .Z(n7_c)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam i2_2_lut_2_lut.init = 16'hdddd;
    FD1S3AY count_wd_delay_i13 (.D(count_wd_delay_31__N_1216[13]), .CK(sys_clk), 
            .Q(count_wd_delay[13])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[14] 151[12])
    defparam count_wd_delay_i13.GSR = "ENABLED";
    FD1S3AY count_wd_delay_i12 (.D(count_wd_delay_31__N_1216[12]), .CK(sys_clk), 
            .Q(count_wd_delay[12])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[14] 151[12])
    defparam count_wd_delay_i12.GSR = "ENABLED";
    FD1S3AY count_wd_delay_i10 (.D(count_wd_delay_31__N_1216[10]), .CK(sys_clk), 
            .Q(count_wd_delay[10])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[14] 151[12])
    defparam count_wd_delay_i10.GSR = "ENABLED";
    FD1S3AY count_wd_delay_i8 (.D(count_wd_delay_31__N_1216[8]), .CK(sys_clk), 
            .Q(count_wd_delay[8])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[14] 151[12])
    defparam count_wd_delay_i8.GSR = "ENABLED";
    FD1S3AY count_wd_delay_i7 (.D(count_wd_delay_31__N_1216[7]), .CK(sys_clk), 
            .Q(count_wd_delay[7])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[14] 151[12])
    defparam count_wd_delay_i7.GSR = "ENABLED";
    FD1S3AY count_wd_delay_i5 (.D(count_wd_delay_31__N_1216[5]), .CK(sys_clk), 
            .Q(count_wd_delay[5])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[14] 151[12])
    defparam count_wd_delay_i5.GSR = "ENABLED";
    FD1S3AY count_wd_delay_i4 (.D(count_wd_delay_31__N_1216[4]), .CK(sys_clk), 
            .Q(count_wd_delay[4])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[14] 151[12])
    defparam count_wd_delay_i4.GSR = "ENABLED";
    FD1S3AY count_wd_delay_i3 (.D(count_wd_delay_31__N_1216[3]), .CK(sys_clk), 
            .Q(count_wd_delay[3])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[14] 151[12])
    defparam count_wd_delay_i3.GSR = "ENABLED";
    FD1S3AY count_wd_delay_i2 (.D(count_wd_delay_31__N_1216[2]), .CK(sys_clk), 
            .Q(count_wd_delay[2])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[14] 151[12])
    defparam count_wd_delay_i2.GSR = "ENABLED";
    LUT4 i1_2_lut_2_lut (.A(\i2c_top_debug[1] ), .B(data_rx_adj_5257[2]), 
         .Z(n4_adj_5238)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam i1_2_lut_2_lut.init = 16'h4444;
    LUT4 n28056_bdd_4_lut_3_lut (.A(\i2c_top_debug[1] ), .B(\i2c_top_debug[3] ), 
         .C(n52298), .Z(n51765)) /* synthesis lut_function=(!(A (B+(C))+!A ((C)+!B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam n28056_bdd_4_lut_3_lut.init = 16'h0606;
    FD1S3AY count_wd_delay_i1 (.D(count_wd_delay_31__N_1216[1]), .CK(sys_clk), 
            .Q(count_wd_delay[1])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[14] 151[12])
    defparam count_wd_delay_i1.GSR = "ENABLED";
    LUT4 i39622_4_lut (.A(\i2c_top_debug[1] ), .B(next_addr_7__N_1168), 
         .C(n52306), .D(\i2c_top_debug[0] ), .Z(data_rx_7__N_1159)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(101[20:44])
    defparam i39622_4_lut.init = 16'h3337;
    LUT4 i2_4_lut_4_lut_4_lut_adj_289 (.A(\i2c_top_debug[1] ), .B(n48025), 
         .C(n7_adj_5239), .D(n52425), .Z(n48963)) /* synthesis lut_function=(!(A (((D)+!C)+!B)+!A ((D)+!B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam i2_4_lut_4_lut_4_lut_adj_289.init = 16'h00c4;
    PFUMX i41683 (.BLUT(n53881), .ALUT(n53882), .C0(\i2c_top_debug[1] ), 
          .Z(n53883));
    LUT4 i39722_2_lut (.A(\i2c_top_debug[5] ), .B(\i2c_top_debug[4] ), .Z(n49650)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i39722_2_lut.init = 16'heeee;
    LUT4 i2c_top_debug_5__I_0_767_Mux_1_i63_4_lut (.A(n31_adj_5205), .B(data_latch), 
         .C(\i2c_top_debug[5] ), .D(n52232), .Z(next_addr_7__N_1160[1])) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i2c_top_debug_5__I_0_767_Mux_1_i63_4_lut.init = 16'h3a0a;
    LUT4 i26167_4_lut_4_lut (.A(n52193), .B(n63), .C(n77[31]), .D(count_wd_delay[31]), 
         .Z(count_wd_delay_31__N_1216[31])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[19:72])
    defparam i26167_4_lut_4_lut.init = 16'h5140;
    LUT4 i2_3_lut_4_lut_4_lut (.A(\i2c_top_debug[0] ), .B(n47760), .C(n52192), 
         .D(byte_rd_left[5]), .Z(n48815)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i2_3_lut_4_lut_4_lut.init = 16'h4440;
    LUT4 n6856_bdd_4_lut_4_lut (.A(\i2c_top_debug[0] ), .B(n52228), .C(\data_reg[3] ), 
         .D(\i2c_top_debug[1] ), .Z(n51918)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam n6856_bdd_4_lut_4_lut.init = 16'h4000;
    LUT4 i2c_top_debug_1__bdd_4_lut_40705_4_lut (.A(\i2c_top_debug[0] ), .B(n52228), 
         .C(n53886), .D(\data_reg[5] ), .Z(n51734)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i2c_top_debug_1__bdd_4_lut_40705_4_lut.init = 16'h4000;
    LUT4 i2c_top_debug_1__bdd_4_lut_4_lut (.A(\i2c_top_debug[0] ), .B(n52228), 
         .C(\i2c_top_debug[2] ), .D(\data_reg[2] ), .Z(n51849)) /* synthesis lut_function=(!(A+!(B (C (D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i2c_top_debug_1__bdd_4_lut_4_lut.init = 16'h4000;
    LUT4 i2c_top_debug_5__I_0_768_Mux_4_i13_4_lut_3_lut (.A(\i2c_top_debug[0] ), 
         .B(data_tx[4]), .C(\i2c_top_debug[1] ), .Z(n37453)) /* synthesis lut_function=(A (C)+!A (B+!(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i2c_top_debug_5__I_0_768_Mux_4_i13_4_lut_3_lut.init = 16'he5e5;
    LUT4 i1_2_lut_adj_290 (.A(\next_i2c_state_4__N_1050[0] ), .B(n66), .Z(n69)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam i1_2_lut_adj_290.init = 16'h8888;
    LUT4 i2_2_lut_adj_291 (.A(write_action), .B(read_action), .Z(n7_adj_5241)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i2_2_lut_adj_291.init = 16'h2222;
    LUT4 mux_464_Mux_0_i31_4_lut_4_lut (.A(\i2c_top_debug[5] ), .B(\i2c_top_debug[2] ), 
         .C(n49518), .D(n49517), .Z(n31_adj_5242)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam mux_464_Mux_0_i31_4_lut_4_lut.init = 16'hf4b0;
    LUT4 i39791_2_lut_rep_480 (.A(\i2c_top_debug[3] ), .B(\i2c_top_debug[2] ), 
         .Z(n52416)) /* synthesis lut_function=((B)+!A) */ ;
    defparam i39791_2_lut_rep_480.init = 16'hdddd;
    LUT4 i39718_2_lut_3_lut (.A(\i2c_top_debug[3] ), .B(\i2c_top_debug[2] ), 
         .C(\i2c_top_debug[5] ), .Z(n49652)) /* synthesis lut_function=((B+(C))+!A) */ ;
    defparam i39718_2_lut_3_lut.init = 16'hfdfd;
    LUT4 n49498_bdd_3_lut_41277_else_4_lut (.A(n52425), .B(\i2c_top_debug[0] ), 
         .C(data_rx_adj_5257[2]), .D(data_rx_adj_5257[5]), .Z(n53881)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam n49498_bdd_3_lut_41277_else_4_lut.init = 16'h0080;
    LUT4 i3_4_lut_4_lut_4_lut (.A(data_rx_adj_5257[6]), .B(n48117), .C(n52262), 
         .D(\i2c_top_debug[4] ), .Z(n49034)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1010[28:70])
    defparam i3_4_lut_4_lut_4_lut.init = 16'h0040;
    LUT4 i26207_4_lut_4_lut (.A(n52193), .B(n63), .C(n77[7]), .D(count_wd_delay[7]), 
         .Z(count_wd_delay_31__N_1216[7])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[19:72])
    defparam i26207_4_lut_4_lut.init = 16'h5140;
    LUT4 i2409_3_lut_4_lut_4_lut (.A(data_rx_adj_5257[6]), .B(data_rx_adj_5257[2]), 
         .C(ack_flag), .D(ack), .Z(n4068)) /* synthesis lut_function=(A (B (C (D)))+!A (C (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1010[28:70])
    defparam i2409_3_lut_4_lut_4_lut.init = 16'hd000;
    FD1P3AX byte_wr_left_6626__i0 (.D(n17[0]), .SP(sys_clk_enable_148), 
            .CK(sys_clk), .Q(byte_wr_left[0]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(750[46:65])
    defparam byte_wr_left_6626__i0.GSR = "ENABLED";
    LUT4 i39703_4_lut (.A(\i2c_top_debug[5] ), .B(\i2c_top_debug[4] ), .C(\i2c_top_debug[3] ), 
         .D(\i2c_top_debug[2] ), .Z(n49672)) /* synthesis lut_function=(A+(B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i39703_4_lut.init = 16'heaaa;
    LUT4 i26651_2_lut_3_lut_4_lut (.A(\i2c_top_debug[1] ), .B(n52306), .C(clear_waiting_ms_N_893), 
         .D(next_addr_7__N_1168), .Z(clear_waiting_ms)) /* synthesis lut_function=(A (C+!(D))+!A ((C+!(D))+!B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i26651_2_lut_3_lut_4_lut.init = 16'hf1ff;
    LUT4 i24418_4_lut_4_lut (.A(n52263), .B(n48845), .C(\i2c_top_debug[2] ), 
         .D(n52301), .Z(n29_adj_5243)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A !(B+(C+(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam i24418_4_lut_4_lut.init = 16'h5f5c;
    LUT4 i3707_4_lut_4_lut (.A(byte_rd_left[5]), .B(n52192), .C(n10_adj_5212), 
         .D(byte_rd_left_5__N_1248[4]), .Z(n7628)) /* synthesis lut_function=(A+(B ((D)+!C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(226[29:50])
    defparam i3707_4_lut_4_lut.init = 16'heeae;
    LUT4 i26983_2_lut (.A(wd_event_active), .B(\i2c_top_debug[5] ), .Z(n37653)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i26983_2_lut.init = 16'heeee;
    LUT4 i26176_4_lut_4_lut (.A(n52193), .B(n63), .C(n77[28]), .D(count_wd_delay[28]), 
         .Z(count_wd_delay_31__N_1216[28])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[19:72])
    defparam i26176_4_lut_4_lut.init = 16'h5140;
    LUT4 i2_2_lut_3_lut (.A(\i2c_top_debug[1] ), .B(n52306), .C(\next_i2c_device_driver_state[4] ), 
         .Z(n7)) /* synthesis lut_function=(A (C)+!A ((C)+!B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i2_2_lut_3_lut.init = 16'hf1f1;
    LUT4 i27241_3_lut_4_lut (.A(\i2c_top_debug[0] ), .B(\i2c_top_debug[2] ), 
         .C(\i2c_top_debug[1] ), .D(n52425), .Z(n37916)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i27241_3_lut_4_lut.init = 16'hff60;
    LUT4 i12566_2_lut_rep_487 (.A(\i2c_top_debug[0] ), .B(\i2c_top_debug[1] ), 
         .Z(n52423)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i12566_2_lut_rep_487.init = 16'h2222;
    LUT4 i26178_4_lut_4_lut (.A(n52193), .B(n63), .C(n77[27]), .D(count_wd_delay[27]), 
         .Z(count_wd_delay_31__N_1216[27])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[19:72])
    defparam i26178_4_lut_4_lut.init = 16'h5140;
    LUT4 i38888_2_lut_rep_488 (.A(\i2c_top_debug[0] ), .B(\i2c_top_debug[1] ), 
         .Z(n52424)) /* synthesis lut_function=(A (B)) */ ;
    defparam i38888_2_lut_rep_488.init = 16'h8888;
    LUT4 i1_2_lut_rep_339_3_lut (.A(\i2c_top_debug[0] ), .B(\i2c_top_debug[1] ), 
         .C(\i2c_top_debug[2] ), .Z(n52275)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_2_lut_rep_339_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_292 (.A(\i2c_top_debug[0] ), .B(\i2c_top_debug[1] ), 
         .C(read_action), .D(\i2c_top_debug[2] ), .Z(n4_adj_5200)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_3_lut_4_lut_adj_292.init = 16'h8000;
    LUT4 i26946_2_lut_rep_293_3_lut_4_lut (.A(\i2c_top_debug[0] ), .B(\i2c_top_debug[1] ), 
         .C(n52425), .D(n53886), .Z(n52229)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i26946_2_lut_rep_293_3_lut_4_lut.init = 16'h8000;
    LUT4 i38599_3_lut_4_lut (.A(n52425), .B(n52275), .C(\i2c_top_debug[3] ), 
         .D(n29_adj_5243), .Z(n49394)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A (C (D))) */ ;
    defparam i38599_3_lut_4_lut.init = 16'hf808;
    LUT4 i26179_4_lut_4_lut (.A(n52193), .B(n63), .C(n77[26]), .D(count_wd_delay[26]), 
         .Z(count_wd_delay_31__N_1216[26])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[19:72])
    defparam i26179_4_lut_4_lut.init = 16'h5140;
    LUT4 ack_I_0_2_lut_rep_489 (.A(ack), .B(ack_flag), .Z(n52425)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam ack_I_0_2_lut_rep_489.init = 16'h8888;
    LUT4 i25806_3_lut_3_lut_4_lut (.A(ack), .B(ack_flag), .C(next_data_latch_N_1505), 
         .D(data_latch), .Z(n12368[0])) /* synthesis lut_function=(!(A (B ((D)+!C)+!B (D))+!A (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam i25806_3_lut_3_lut_4_lut.init = 16'h00f7;
    LUT4 i1_2_lut_3_lut_3_lut_4_lut (.A(ack), .B(ack_flag), .C(n52455), 
         .D(\i2c_top_debug[0] ), .Z(n27301)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam i1_2_lut_3_lut_3_lut_4_lut.init = 16'h7000;
    LUT4 i38706_3_lut_4_lut (.A(ack), .B(ack_flag), .C(\i2c_top_debug[3] ), 
         .D(count_us[11]), .Z(n49501)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam i38706_3_lut_4_lut.init = 16'h8f80;
    LUT4 i27462_2_lut_3_lut_4_lut (.A(ack), .B(ack_flag), .C(\i2c_top_debug[1] ), 
         .D(\i2c_top_debug[0] ), .Z(n38161)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam i27462_2_lut_3_lut_4_lut.init = 16'h0800;
    LUT4 i2_3_lut_4_lut_adj_293 (.A(ack), .B(ack_flag), .C(n47760), .D(\i2c_top_debug[0] ), 
         .Z(n48814)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam i2_3_lut_4_lut_adj_293.init = 16'h8000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_294 (.A(ack), .B(ack_flag), .C(n52459), 
         .D(data_rx_adj_5257[2]), .Z(n4_adj_5210)) /* synthesis lut_function=(((C+!(D))+!B)+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam i1_2_lut_3_lut_4_lut_adj_294.init = 16'hf7ff;
    LUT4 i3_3_lut_3_lut_4_lut (.A(ack), .B(ack_flag), .C(n52452), .D(n52436), 
         .Z(n49064)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A (C+!(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam i3_3_lut_3_lut_4_lut.init = 16'h0700;
    LUT4 i39771_2_lut_3_lut (.A(ack), .B(ack_flag), .C(\i2c_top_debug[0] ), 
         .Z(n34018)) /* synthesis lut_function=(!(A (B+(C))+!A (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam i39771_2_lut_3_lut.init = 16'h0707;
    LUT4 i1_2_lut_rep_327_3_lut_4_lut (.A(ack), .B(ack_flag), .C(\i2c_top_debug[1] ), 
         .D(\i2c_top_debug[0] ), .Z(n52263)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam i1_2_lut_rep_327_3_lut_4_lut.init = 16'h8000;
    LUT4 i26796_3_lut_3_lut_4_lut (.A(ack), .B(ack_flag), .C(n26115), 
         .D(\i2c_top_debug[3] ), .Z(n15_adj_5206)) /* synthesis lut_function=(!(A (B+!(C+(D)))+!A !(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam i26796_3_lut_3_lut_4_lut.init = 16'h7770;
    LUT4 i1_2_lut_2_lut_3_lut (.A(ack), .B(ack_flag), .C(data_rx_adj_5257[6]), 
         .Z(n48)) /* synthesis lut_function=(((C)+!B)+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam i1_2_lut_2_lut_3_lut.init = 16'hf7f7;
    LUT4 i11546_4_lut_3_lut_4_lut (.A(ack), .B(ack_flag), .C(\i2c_top_debug[0] ), 
         .D(n4_adj_5238), .Z(n21941)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A !(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam i11546_4_lut_3_lut_4_lut.init = 16'h7870;
    LUT4 i9138_3_lut_4_lut (.A(ack), .B(ack_flag), .C(n52277), .D(data_latch), 
         .Z(n18960)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam i9138_3_lut_4_lut.init = 16'h707f;
    LUT4 n6856_bdd_2_lut_2_lut_3_lut_4_lut (.A(ack), .B(ack_flag), .C(\i2c_top_debug[1] ), 
         .D(\i2c_top_debug[0] ), .Z(n51917)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A !(C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam n6856_bdd_2_lut_2_lut_3_lut_4_lut.init = 16'h7000;
    LUT4 i1_2_lut_3_lut_4_lut_adj_295 (.A(ack), .B(ack_flag), .C(n52459), 
         .D(\i2c_top_debug[0] ), .Z(n4_adj_5203)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam i1_2_lut_3_lut_4_lut_adj_295.init = 16'h0080;
    LUT4 i1_2_lut_3_lut_4_lut_adj_296 (.A(ack), .B(ack_flag), .C(n45033), 
         .D(data_latch), .Z(n2486[5])) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam i1_2_lut_3_lut_4_lut_adj_296.init = 16'h0080;
    LUT4 i2c_top_debug_1__bdd_2_lut_3_lut_4_lut (.A(ack), .B(ack_flag), 
         .C(\i2c_top_debug[1] ), .D(\i2c_top_debug[0] ), .Z(n50985)) /* synthesis lut_function=(!(A (B (C (D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam i2c_top_debug_1__bdd_2_lut_3_lut_4_lut.init = 16'h7fff;
    LUT4 i1_2_lut_rep_298_3_lut_4_lut (.A(ack), .B(ack_flag), .C(n52431), 
         .D(\i2c_top_debug[0] ), .Z(n52234)) /* synthesis lut_function=(!(((C+!(D))+!B)+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam i1_2_lut_rep_298_3_lut_4_lut.init = 16'h0800;
    LUT4 i1_2_lut_rep_362_3_lut (.A(ack), .B(ack_flag), .C(\i2c_top_debug[0] ), 
         .Z(n52298)) /* synthesis lut_function=(A (B+!(C))+!A !(C)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam i1_2_lut_rep_362_3_lut.init = 16'h8f8f;
    LUT4 i1_2_lut_rep_357_3_lut (.A(ack), .B(ack_flag), .C(\i2c_top_debug[0] ), 
         .Z(n52293)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam i1_2_lut_rep_357_3_lut.init = 16'h8080;
    LUT4 i38707_3_lut_4_lut (.A(ack), .B(ack_flag), .C(\i2c_top_debug[3] ), 
         .D(go), .Z(n49502)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam i38707_3_lut_4_lut.init = 16'h8f80;
    LUT4 i1_2_lut_3_lut_4_lut_adj_297 (.A(ack), .B(ack_flag), .C(\i2c_top_debug[1] ), 
         .D(\i2c_top_debug[0] ), .Z(n28051)) /* synthesis lut_function=(A (B+(C+!(D)))+!A (C+!(D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam i1_2_lut_3_lut_4_lut_adj_297.init = 16'hf8ff;
    LUT4 i27293_1_lut_2_lut_3_lut_4_lut (.A(ack), .B(ack_flag), .C(n1516), 
         .D(\i2c_top_debug[0] ), .Z(n24)) /* synthesis lut_function=(!(A (B (C (D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam i27293_1_lut_2_lut_3_lut_4_lut.init = 16'h7fff;
    LUT4 i38710_3_lut_3_lut_4_lut (.A(ack), .B(ack_flag), .C(n12358[0]), 
         .D(\i2c_top_debug[0] ), .Z(n49505)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam i38710_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 i39638_2_lut_rep_363_3_lut (.A(ack), .B(ack_flag), .C(data_rx_adj_5257[2]), 
         .Z(n52299)) /* synthesis lut_function=(!(A (B (C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam i39638_2_lut_rep_363_3_lut.init = 16'h7f7f;
    LUT4 i33212_3_lut_3_lut_4_lut (.A(ack), .B(ack_flag), .C(n47361), 
         .D(\i2c_top_debug[3] ), .Z(n43988)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam i33212_3_lut_3_lut_4_lut.init = 16'h77f0;
    LUT4 i1_2_lut_rep_264_3_lut_3_lut_3_lut_4_lut (.A(ack), .B(ack_flag), 
         .C(n52455), .D(\i2c_top_debug[0] ), .Z(n52200)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam i1_2_lut_rep_264_3_lut_3_lut_3_lut_4_lut.init = 16'h0070;
    PFUMX mux_464_Mux_0_i63 (.BLUT(n49461), .ALUT(n31_adj_5242), .C0(n49529), 
          .Z(next_i2c_cmd_state_5__N_1479[0])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;
    LUT4 i26937_2_lut_rep_305_3_lut_4_lut (.A(ack), .B(ack_flag), .C(n1516), 
         .D(\i2c_top_debug[0] ), .Z(n52241)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam i26937_2_lut_rep_305_3_lut_4_lut.init = 16'h8000;
    LUT4 i38709_3_lut_4_lut_3_lut_4_lut (.A(ack), .B(ack_flag), .C(n52466), 
         .D(\i2c_top_debug[0] ), .Z(n49504)) /* synthesis lut_function=(A (B (C+!(D))+!B (D))+!A (D)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam i38709_3_lut_4_lut_3_lut_4_lut.init = 16'hf788;
    LUT4 i26775_2_lut_2_lut_3_lut_4_lut (.A(ack), .B(ack_flag), .C(\i2c_top_debug[1] ), 
         .D(\i2c_top_debug[0] ), .Z(n7_adj_5245)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A (C+!(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam i26775_2_lut_2_lut_3_lut_4_lut.init = 16'h0700;
    LUT4 clear_waiting_us_N_1214_bdd_4_lut_40430_2_lut_3_lut (.A(ack), .B(ack_flag), 
         .C(\i2c_top_debug[0] ), .Z(n51194)) /* synthesis lut_function=(!(A (B+!(C))+!A !(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam clear_waiting_us_N_1214_bdd_4_lut_40430_2_lut_3_lut.init = 16'h7070;
    LUT4 i1_2_lut_rep_326_3_lut (.A(ack), .B(ack_flag), .C(\i2c_top_debug[0] ), 
         .Z(n52262)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam i1_2_lut_rep_326_3_lut.init = 16'h0808;
    PFUMX i40192 (.BLUT(n51037), .ALUT(n51036), .C0(\i2c_top_debug[4] ), 
          .Z(n51038));
    LUT4 i26181_4_lut_4_lut (.A(n52193), .B(n63), .C(n77[25]), .D(count_wd_delay[25]), 
         .Z(count_wd_delay_31__N_1216[25])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[19:72])
    defparam i26181_4_lut_4_lut.init = 16'h5140;
    LUT4 next_data_tx_7__N_1439_4__bdd_2_lut_2_lut_3_lut_4_lut (.A(ack), .B(ack_flag), 
         .C(\i2c_top_debug[1] ), .D(\i2c_top_debug[0] ), .Z(n52026)) /* synthesis lut_function=(!(A (B+!((D)+!C))+!A !((D)+!C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam next_data_tx_7__N_1439_4__bdd_2_lut_2_lut_3_lut_4_lut.init = 16'h7707;
    LUT4 i3_3_lut_3_lut_4_lut_adj_298 (.A(ack), .B(ack_flag), .C(\i2c_top_debug[0] ), 
         .D(n53886), .Z(n8_adj_5246)) /* synthesis lut_function=(((C+(D))+!B)+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam i3_3_lut_3_lut_4_lut_adj_298.init = 16'hfff7;
    LUT4 i39911_2_lut_rep_323_3_lut_4_lut (.A(ack), .B(ack_flag), .C(\i2c_top_debug[1] ), 
         .D(\i2c_top_debug[0] ), .Z(n52259)) /* synthesis lut_function=(!(A (B+((D)+!C))+!A ((D)+!C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam i39911_2_lut_rep_323_3_lut_4_lut.init = 16'h0070;
    LUT4 i22311_3_lut_4_lut (.A(ack), .B(ack_flag), .C(\i2c_top_debug[3] ), 
         .D(count_us_11__N_1299), .Z(n5)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam i22311_3_lut_4_lut.init = 16'h8f80;
    LUT4 i6_1_lut_rep_364_2_lut (.A(ack), .B(ack_flag), .Z(n52300)) /* synthesis lut_function=(!(A (B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam i6_1_lut_rep_364_2_lut.init = 16'h7777;
    LUT4 i38623_4_lut_4_lut (.A(n52229), .B(n8_adj_5246), .C(\i2c_top_debug[3] ), 
         .D(n7_c), .Z(n49418)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A !(B+(C+(D))))) */ ;
    defparam i38623_4_lut_4_lut.init = 16'h5f5c;
    LUT4 i38598_4_lut_4_lut (.A(n52229), .B(n8_adj_5247), .C(\i2c_top_debug[3] ), 
         .D(n7_adj_5241), .Z(n49393)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A !(B (C+(D))+!B (C)))) */ ;
    defparam i38598_4_lut_4_lut.init = 16'h5c50;
    L6MUX21 i38665 (.D0(n25_adj_5218), .D1(n49506), .SD(\i2c_top_debug[2] ), 
            .Z(n49460));
    LUT4 i22353_3_lut_4_lut_3_lut_4_lut (.A(ack), .B(ack_flag), .C(data_rx_adj_5257[2]), 
         .D(\i2c_top_debug[1] ), .Z(n33015)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A !(D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam i22353_3_lut_4_lut_3_lut_4_lut.init = 16'h7780;
    LUT4 mux_464_Mux_0_i24_3_lut_4_lut (.A(ack), .B(ack_flag), .C(\i2c_top_debug[0] ), 
         .D(n1516), .Z(n24_adj_5217)) /* synthesis lut_function=(!(A (B (C (D))+!B !(C))+!A !(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam mux_464_Mux_0_i24_3_lut_4_lut.init = 16'h78f8;
    LUT4 i27526_2_lut_3_lut_4_lut (.A(ack), .B(ack_flag), .C(\i2c_top_debug[1] ), 
         .D(\i2c_top_debug[0] ), .Z(n38227)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A !(C+!(D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(1003[25:66])
    defparam i27526_2_lut_3_lut_4_lut.init = 16'h8f88;
    PFUMX i38711 (.BLUT(n49504), .ALUT(n49505), .C0(\i2c_top_debug[1] ), 
          .Z(n49506));
    PFUMX i40823 (.BLUT(n52028), .ALUT(n52024), .C0(n49672), .Z(next_addr_7__N_1160[2]));
    PFUMX i40821 (.BLUT(n52026), .ALUT(n52025), .C0(n52432), .Z(n52027));
    L6MUX21 mux_464_Mux_2_i63 (.D0(n49389), .D1(n31_adj_5248), .SD(n49650), 
            .Z(next_i2c_cmd_state_5__N_1479[2])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;
    LUT4 i3_4_lut_4_lut (.A(\i2c_top_debug[4] ), .B(n37653), .C(n52291), 
         .D(n48025), .Z(n66)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(267[14] 1038[12])
    defparam i3_4_lut_4_lut.init = 16'h1000;
    PFUMX i34257 (.BLUT(n48815), .ALUT(n48112), .C0(\i2c_top_debug[5] ), 
          .Z(n45033));
    LUT4 n52027_bdd_3_lut_3_lut (.A(\i2c_top_debug[4] ), .B(n52539), .C(n52027), 
         .Z(n52028)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(267[14] 1038[12])
    defparam n52027_bdd_3_lut_3_lut.init = 16'he4e4;
    LUT4 i1_2_lut_adj_299 (.A(count_us_11__N_1287[11]), .B(count_us_11__N_1299), 
         .Z(n26[11])) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(128[14] 131[34])
    defparam i1_2_lut_adj_299.init = 16'hbbbb;
    LUT4 i2_3_lut_3_lut_3_lut (.A(\i2c_top_debug[2] ), .B(\i2c_top_debug[3] ), 
         .C(\i2c_top_debug[4] ), .Z(n48712)) /* synthesis lut_function=((B+!(C))+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(267[14] 1038[12])
    defparam i2_3_lut_3_lut_3_lut.init = 16'hdfdf;
    PFUMX i38594 (.BLUT(n49387), .ALUT(n49388), .C0(\i2c_top_debug[3] ), 
          .Z(n49389));
    LUT4 i1_2_lut_3_lut_4_lut_4_lut (.A(\i2c_top_debug[2] ), .B(n52464), 
         .C(next_data_latch_N_1505), .D(n52423), .Z(n48112)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(267[14] 1038[12])
    defparam i1_2_lut_3_lut_4_lut_4_lut.init = 16'h1000;
    CCU2D sub_10_add_2_13 (.A0(count_us[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n43947), .S0(count_us_11__N_1287[11]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(129[25:42])
    defparam sub_10_add_2_13.INIT0 = 16'h5555;
    defparam sub_10_add_2_13.INIT1 = 16'h0000;
    defparam sub_10_add_2_13.INJECT1_0 = "NO";
    defparam sub_10_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_11 (.A0(count_us[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_us[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43946), .COUT(n43947), .S0(count_us_11__N_1287[9]), 
          .S1(count_us_11__N_1287[10]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(129[25:42])
    defparam sub_10_add_2_11.INIT0 = 16'h5555;
    defparam sub_10_add_2_11.INIT1 = 16'h5555;
    defparam sub_10_add_2_11.INJECT1_0 = "NO";
    defparam sub_10_add_2_11.INJECT1_1 = "NO";
    LUT4 i1_2_lut_rep_296_3_lut_4_lut_4_lut (.A(n53886), .B(n52464), .C(\i2c_top_debug[1] ), 
         .D(\i2c_top_debug[0] ), .Z(n52232)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(267[14] 1038[12])
    defparam i1_2_lut_rep_296_3_lut_4_lut_4_lut.init = 16'h0100;
    LUT4 i27126_3_lut_4_lut_4_lut (.A(\i2c_top_debug[2] ), .B(n52436), .C(ack_flag), 
         .D(ack), .Z(n29_adj_5249)) /* synthesis lut_function=(!((B+(C (D)))+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(267[14] 1038[12])
    defparam i27126_3_lut_4_lut_4_lut.init = 16'h0222;
    LUT4 i1_2_lut_rep_337_3_lut_3_lut (.A(n53886), .B(\i2c_top_debug[1] ), 
         .C(\i2c_top_debug[0] ), .Z(n52273)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(267[14] 1038[12])
    defparam i1_2_lut_rep_337_3_lut_3_lut.init = 16'h1010;
    LUT4 i26885_2_lut_rep_294_3_lut_3_lut_4_lut_4_lut (.A(n53886), .B(n52425), 
         .C(\i2c_top_debug[1] ), .D(\i2c_top_debug[0] ), .Z(n52230)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(267[14] 1038[12])
    defparam i26885_2_lut_rep_294_3_lut_3_lut_4_lut_4_lut.init = 16'h0100;
    LUT4 i3_2_lut_3_lut_4_lut (.A(\i2c_top_debug[2] ), .B(\i2c_top_debug[1] ), 
         .C(n4068), .D(\i2c_top_debug[0] ), .Z(n8_adj_5247)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(267[14] 1038[12])
    defparam i3_2_lut_3_lut_4_lut.init = 16'h8000;
    LUT4 i1_2_lut_rep_353_3_lut (.A(n53886), .B(\i2c_top_debug[1] ), .C(\i2c_top_debug[0] ), 
         .Z(n52289)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(267[14] 1038[12])
    defparam i1_2_lut_rep_353_3_lut.init = 16'h8080;
    LUT4 i1_2_lut_rep_495 (.A(n53886), .B(\i2c_top_debug[1] ), .Z(n52431)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(267[14] 1038[12])
    defparam i1_2_lut_rep_495.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_adj_300 (.A(n53886), .B(\i2c_top_debug[1] ), .C(\i2c_top_debug[3] ), 
         .Z(n44475)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(267[14] 1038[12])
    defparam i1_2_lut_3_lut_adj_300.init = 16'h1010;
    LUT4 i3452_1_lut_rep_496 (.A(\i2c_top_debug[3] ), .Z(n52432)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam i3452_1_lut_rep_496.init = 16'h5555;
    LUT4 i27345_2_lut_4_lut_4_lut_4_lut (.A(\i2c_top_debug[3] ), .B(n52316), 
         .C(data_latch), .D(\i2c_top_debug[2] ), .Z(n30_adj_5204)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam i27345_2_lut_4_lut_4_lut_4_lut.init = 16'h0200;
    LUT4 i39177_3_lut_4_lut_4_lut (.A(\i2c_top_debug[3] ), .B(n7_adj_5245), 
         .C(data_tx[7]), .D(n52259), .Z(n14_adj_5251)) /* synthesis lut_function=(A (C (D))+!A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam i39177_3_lut_4_lut_4_lut.init = 16'he444;
    PFUMX i40762 (.BLUT(n51923), .ALUT(n53875), .C0(\i2c_top_debug[4] ), 
          .Z(n51924));
    LUT4 i2_3_lut_rep_341_4_lut_4_lut_4_lut (.A(\i2c_top_debug[3] ), .B(\i2c_top_debug[0] ), 
         .C(\i2c_top_debug[1] ), .D(\i2c_top_debug[2] ), .Z(n52277)) /* synthesis lut_function=((B+!(C (D)))+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam i2_3_lut_rep_341_4_lut_4_lut_4_lut.init = 16'hdfff;
    LUT4 gnd_bdd_2_lut_40734_3_lut_3_lut (.A(\i2c_top_debug[3] ), .B(\i2c_top_debug[1] ), 
         .C(n51849), .Z(n51851)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam gnd_bdd_2_lut_40734_3_lut_3_lut.init = 16'h4040;
    LUT4 i1_2_lut_rep_355_2_lut (.A(\i2c_top_debug[3] ), .B(\i2c_top_debug[1] ), 
         .Z(n52291)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam i1_2_lut_rep_355_2_lut.init = 16'h4444;
    LUT4 i2_3_lut_4_lut_4_lut_adj_301 (.A(\i2c_top_debug[3] ), .B(\i2c_top_debug[2] ), 
         .C(\i2c_top_debug[1] ), .D(\i2c_top_debug[0] ), .Z(n48829)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam i2_3_lut_4_lut_4_lut_adj_301.init = 16'h0400;
    LUT4 i2c_top_debug_5__I_0_768_Mux_1_i14_4_lut_4_lut (.A(\i2c_top_debug[3] ), 
         .B(n52259), .C(n52230), .D(data_tx[1]), .Z(n14)) /* synthesis lut_function=(A (B (D))+!A (C)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam i2c_top_debug_5__I_0_768_Mux_1_i14_4_lut_4_lut.init = 16'hd850;
    PFUMX i40759 (.BLUT(n51921), .ALUT(n51759), .C0(\i2c_top_debug[2] ), 
          .Z(n51922));
    LUT4 i1_3_lut_4_lut_4_lut (.A(\i2c_top_debug[3] ), .B(n53), .C(ack_flag), 
         .D(ack), .Z(n32988)) /* synthesis lut_function=(A (B (C (D)))+!A (C (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam i1_3_lut_4_lut_4_lut.init = 16'hd000;
    LUT4 i1_2_lut_3_lut_3_lut_3_lut (.A(\i2c_top_debug[3] ), .B(\i2c_top_debug[1] ), 
         .C(\i2c_top_debug[2] ), .Z(n48117)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam i1_2_lut_3_lut_3_lut_3_lut.init = 16'h0404;
    LUT4 i2c_top_debug_5__I_0_768_Mux_4_i14_4_lut_4_lut_4_lut_4_lut (.A(\i2c_top_debug[3] ), 
         .B(n52273), .C(n37453), .D(n52425), .Z(n14_adj_5253)) /* synthesis lut_function=(!(A ((D)+!C)+!A ((D)+!B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam i2c_top_debug_5__I_0_768_Mux_4_i14_4_lut_4_lut_4_lut_4_lut.init = 16'h00e4;
    LUT4 i63_4_lut_4_lut (.A(\i2c_top_debug[3] ), .B(n51194), .C(\i2c_top_debug[4] ), 
         .D(n28051), .Z(n33)) /* synthesis lut_function=(!(A (D)+!A !(B (C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam i63_4_lut_4_lut.init = 16'h40ea;
    FD1S3IX i2c_cmd_state__i3_rep_532 (.D(next_i2c_cmd_state_5__N_1479[2]), 
            .CK(sys_clk), .CD(wd_event_active), .Q(n53886)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam i2c_cmd_state__i3_rep_532.GSR = "ENABLED";
    LUT4 i22307_4_lut_4_lut (.A(\i2c_top_debug[3] ), .B(n52425), .C(\i2c_top_debug[1] ), 
         .D(data_rx_adj_5257[2]), .Z(n32969)) /* synthesis lut_function=(A (B ((D)+!C))+!A (B+!(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam i22307_4_lut_4_lut.init = 16'hcd4d;
    CCU2D sub_10_add_2_9 (.A0(count_us[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_us[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43945), .COUT(n43946), .S0(count_us_11__N_1287[7]), 
          .S1(count_us_11__N_1287[8]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(129[25:42])
    defparam sub_10_add_2_9.INIT0 = 16'h5555;
    defparam sub_10_add_2_9.INIT1 = 16'h5555;
    defparam sub_10_add_2_9.INJECT1_0 = "NO";
    defparam sub_10_add_2_9.INJECT1_1 = "NO";
    LUT4 i8370_2_lut_rep_500 (.A(\i2c_top_debug[0] ), .B(\i2c_top_debug[1] ), 
         .Z(n52436)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i8370_2_lut_rep_500.init = 16'h6666;
    PFUMX i38708 (.BLUT(n49501), .ALUT(n49502), .C0(\i2c_top_debug[1] ), 
          .Z(n49503));
    CCU2D sub_10_add_2_7 (.A0(count_us[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_us[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43944), .COUT(n43945), .S0(count_us_11__N_1287[5]), 
          .S1(count_us_11__N_1287[6]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(129[25:42])
    defparam sub_10_add_2_7.INIT0 = 16'h5555;
    defparam sub_10_add_2_7.INIT1 = 16'h5555;
    defparam sub_10_add_2_7.INJECT1_0 = "NO";
    defparam sub_10_add_2_7.INJECT1_1 = "NO";
    LUT4 i1_2_lut_3_lut_4_lut_adj_302 (.A(byte_rd_left[2]), .B(n52286), 
         .C(byte_rd_left[4]), .D(byte_rd_left[3]), .Z(byte_rd_left_5__N_1248[4])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)+!C !(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(226[29:50])
    defparam i1_2_lut_3_lut_4_lut_adj_302.init = 16'hf0e1;
    LUT4 i7675_2_lut_rep_256_3_lut_4_lut (.A(byte_rd_left[2]), .B(n52286), 
         .C(byte_rd_left[4]), .D(byte_rd_left[3]), .Z(n52192)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(226[29:50])
    defparam i7675_2_lut_rep_256_3_lut_4_lut.init = 16'hfffe;
    PFUMX i38721 (.BLUT(n32969), .ALUT(n8), .C0(\i2c_top_debug[0] ), .Z(n49516));
    LUT4 i1_2_lut_adj_303 (.A(count_us_11__N_1287[10]), .B(count_us_11__N_1299), 
         .Z(n26[10])) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(128[14] 131[34])
    defparam i1_2_lut_adj_303.init = 16'hbbbb;
    LUT4 i39823_4_lut (.A(count_us[11]), .B(n49222), .C(n49216), .D(count_us[6]), 
         .Z(count_us_11__N_1299)) /* synthesis lut_function=(!(A (B (C (D))))) */ ;
    defparam i39823_4_lut.init = 16'h7fff;
    CCU2D sub_10_add_2_5 (.A0(count_us[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_us[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43943), .COUT(n43944), .S0(count_us_11__N_1287[3]), 
          .S1(count_us_11__N_1287[4]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(129[25:42])
    defparam sub_10_add_2_5.INIT0 = 16'h5555;
    defparam sub_10_add_2_5.INIT1 = 16'h5555;
    defparam sub_10_add_2_5.INJECT1_0 = "NO";
    defparam sub_10_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_3 (.A0(count_us[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_us[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43942), .COUT(n43943), .S0(count_us_11__N_1287[1]), 
          .S1(count_us_11__N_1287[2]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(129[25:42])
    defparam sub_10_add_2_3.INIT0 = 16'h5555;
    defparam sub_10_add_2_3.INIT1 = 16'h5555;
    defparam sub_10_add_2_3.INJECT1_0 = "NO";
    defparam sub_10_add_2_3.INJECT1_1 = "NO";
    LUT4 i1_3_lut (.A(count_us[10]), .B(count_us[0]), .C(count_us[9]), 
         .Z(n49222)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i1_3_lut.init = 16'h8080;
    LUT4 i2_3_lut_4_lut_adj_304 (.A(\i2c_top_debug[1] ), .B(n52200), .C(\data_reg[6] ), 
         .D(\i2c_top_debug[4] ), .Z(n48756)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i2_3_lut_4_lut_adj_304.init = 16'h8000;
    LUT4 i1_4_lut_adj_305 (.A(count_us[8]), .B(n49212), .C(count_us[4]), 
         .D(count_us[5]), .Z(n49216)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_305.init = 16'h8000;
    LUT4 i1_4_lut_adj_306 (.A(count_us[7]), .B(count_us[1]), .C(count_us[2]), 
         .D(count_us[3]), .Z(n49212)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_306.init = 16'h8000;
    LUT4 i19928_3_lut (.A(n30599), .B(n30598), .C(n30594), .Z(count_us[10])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(128[14] 131[34])
    defparam i19928_3_lut.init = 16'hcaca;
    LUT4 i19940_3_lut (.A(n30611), .B(n30610), .C(n30594), .Z(count_us[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(128[14] 131[34])
    defparam i19940_3_lut.init = 16'hcaca;
    LUT4 i19931_3_lut (.A(n30602), .B(n30601), .C(n30594), .Z(count_us[9])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(128[14] 131[34])
    defparam i19931_3_lut.init = 16'hcaca;
    LUT4 i19934_3_lut (.A(n30605), .B(n30604), .C(n30594), .Z(count_us[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(128[14] 131[34])
    defparam i19934_3_lut.init = 16'hcaca;
    CCU2D sub_10_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count_us[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n43942), .S1(count_us_11__N_1287[0]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(129[25:42])
    defparam sub_10_add_2_1.INIT0 = 16'hF000;
    defparam sub_10_add_2_1.INIT1 = 16'h5555;
    defparam sub_10_add_2_1.INJECT1_0 = "NO";
    defparam sub_10_add_2_1.INJECT1_1 = "NO";
    PFUMX i40719 (.BLUT(n51855), .ALUT(n51851), .C0(\i2c_top_debug[4] ), 
          .Z(n51856));
    LUT4 i19925_3_lut (.A(n30596), .B(n30595), .C(n30594), .Z(count_us[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(128[14] 131[34])
    defparam i19925_3_lut.init = 16'hcaca;
    LUT4 i38570_2_lut_3_lut_4_lut (.A(\i2c_top_debug[1] ), .B(n52306), .C(n7246), 
         .D(next_addr_7__N_1168), .Z(n49365)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i38570_2_lut_3_lut_4_lut.init = 16'he000;
    PFUMX i40716 (.BLUT(n51853), .ALUT(n51852), .C0(n53886), .Z(n51854));
    LUT4 i19937_3_lut (.A(n30608), .B(n30607), .C(n30594), .Z(count_us[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(128[14] 131[34])
    defparam i19937_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_307 (.A(count_us_11__N_1287[9]), .B(count_us_11__N_1299), 
         .Z(n26[9])) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(128[14] 131[34])
    defparam i1_2_lut_adj_307.init = 16'hbbbb;
    LUT4 i1_2_lut_adj_308 (.A(count_us_11__N_1299), .B(count_us_11__N_1287[8]), 
         .Z(n26[8])) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(128[14] 131[34])
    defparam i1_2_lut_adj_308.init = 16'hdddd;
    LUT4 i1_2_lut_adj_309 (.A(count_us_11__N_1299), .B(count_us_11__N_1287[6]), 
         .Z(n26[6])) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(128[14] 131[34])
    defparam i1_2_lut_adj_309.init = 16'hdddd;
    LUT4 i39625_2_lut (.A(clear_waiting_us), .B(resetn), .Z(count_us_11__N_1209)) /* synthesis lut_function=(!(A (B))) */ ;
    defparam i39625_2_lut.init = 16'h7777;
    LUT4 count_us_i1_i1_3_lut (.A(count_us[0]), .B(count_us_11__N_1287[0]), 
         .C(count_us_11__N_1299), .Z(n26[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(128[14] 131[34])
    defparam count_us_i1_i1_3_lut.init = 16'hcaca;
    L6MUX21 i38645 (.D0(n49438), .D1(n49439), .SD(\i2c_top_debug[4] ), 
            .Z(n49440));
    PFUMX i40160 (.BLUT(n50986), .ALUT(n50985), .C0(\i2c_top_debug[2] ), 
          .Z(n50987));
    LUT4 i26192_4_lut_4_lut (.A(n52193), .B(n63), .C(n77[12]), .D(count_wd_delay[12]), 
         .Z(count_wd_delay_31__N_1216[12])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[19:72])
    defparam i26192_4_lut_4_lut.init = 16'h5140;
    PFUMX byte_wr_left_6626_mux_6_i2 (.BLUT(n48108), .ALUT(n2[1]), .C0(n6849), 
          .Z(n17[1]));
    L6MUX21 i38597 (.D0(n49390), .D1(n49391), .SD(\i2c_top_debug[4] ), 
            .Z(n49392));
    PFUMX i38600 (.BLUT(n49393), .ALUT(n49394), .C0(\i2c_top_debug[4] ), 
          .Z(n49395));
    LUT4 i24_4_lut_adj_310 (.A(\data_reg[0] ), .B(n48496), .C(\next_i2c_device_driver_state[4] ), 
         .D(n52450), .Z(n10_adj_5208)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(129[9:37])
    defparam i24_4_lut_adj_310.init = 16'hcfca;
    CCU2D sub_31_add_2_33 (.A0(count_wd_delay[31]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n43925), .S0(n77[31]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(145[31:54])
    defparam sub_31_add_2_33.INIT0 = 16'h5555;
    defparam sub_31_add_2_33.INIT1 = 16'h0000;
    defparam sub_31_add_2_33.INJECT1_0 = "NO";
    defparam sub_31_add_2_33.INJECT1_1 = "NO";
    LUT4 n51734_bdd_4_lut (.A(n51734), .B(\i2c_top_debug[1] ), .C(n29_adj_5249), 
         .D(\i2c_top_debug[3] ), .Z(n53872)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)))+!A (C (D))) */ ;
    defparam n51734_bdd_4_lut.init = 16'hf088;
    CCU2D sub_31_add_2_31 (.A0(count_wd_delay[29]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_wd_delay[30]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43924), .COUT(n43925), .S0(n77[29]), .S1(n77[30]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(145[31:54])
    defparam sub_31_add_2_31.INIT0 = 16'h5555;
    defparam sub_31_add_2_31.INIT1 = 16'h5555;
    defparam sub_31_add_2_31.INJECT1_0 = "NO";
    defparam sub_31_add_2_31.INJECT1_1 = "NO";
    CCU2D sub_31_add_2_29 (.A0(count_wd_delay[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_wd_delay[28]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43923), .COUT(n43924), .S0(n77[27]), .S1(n77[28]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(145[31:54])
    defparam sub_31_add_2_29.INIT0 = 16'h5555;
    defparam sub_31_add_2_29.INIT1 = 16'h5555;
    defparam sub_31_add_2_29.INJECT1_0 = "NO";
    defparam sub_31_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_31_add_2_27 (.A0(count_wd_delay[25]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_wd_delay[26]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43922), .COUT(n43923), .S0(n77[25]), .S1(n77[26]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(145[31:54])
    defparam sub_31_add_2_27.INIT0 = 16'h5555;
    defparam sub_31_add_2_27.INIT1 = 16'h5555;
    defparam sub_31_add_2_27.INJECT1_0 = "NO";
    defparam sub_31_add_2_27.INJECT1_1 = "NO";
    L6MUX21 i38722 (.D0(n49503), .D1(n43989), .SD(\i2c_top_debug[0] ), 
            .Z(n49517));
    PFUMX i40657 (.BLUT(n51765), .ALUT(n51764), .C0(n53886), .Z(n51766));
    CCU2D sub_31_add_2_25 (.A0(count_wd_delay[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_wd_delay[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43921), .COUT(n43922), .S0(n77[23]), .S1(n77[24]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(145[31:54])
    defparam sub_31_add_2_25.INIT0 = 16'h5555;
    defparam sub_31_add_2_25.INIT1 = 16'h5555;
    defparam sub_31_add_2_25.INJECT1_0 = "NO";
    defparam sub_31_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_31_add_2_23 (.A0(count_wd_delay[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_wd_delay[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43920), .COUT(n43921), .S0(count_wd_delay_31__N_1300[21]), 
          .S1(n77[22]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(145[31:54])
    defparam sub_31_add_2_23.INIT0 = 16'h5555;
    defparam sub_31_add_2_23.INIT1 = 16'h5555;
    defparam sub_31_add_2_23.INJECT1_0 = "NO";
    defparam sub_31_add_2_23.INJECT1_1 = "NO";
    PFUMX i38644 (.BLUT(n46343), .ALUT(n29_adj_5214), .C0(\i2c_top_debug[3] ), 
          .Z(n49439));
    LUT4 n51536_bdd_4_lut_41280 (.A(n32), .B(\i2c_top_debug[3] ), .C(\i2c_top_debug[0] ), 
         .D(\i2c_top_debug[1] ), .Z(n53175)) /* synthesis lut_function=(!(A (B+(C (D)))+!A (B+(C+!(D))))) */ ;
    defparam n51536_bdd_4_lut_41280.init = 16'h0322;
    LUT4 i26182_4_lut_4_lut (.A(n52193), .B(n63), .C(n77[24]), .D(count_wd_delay[24]), 
         .Z(count_wd_delay_31__N_1216[24])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[19:72])
    defparam i26182_4_lut_4_lut.init = 16'h5140;
    CCU2D sub_31_add_2_21 (.A0(count_wd_delay[19]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_wd_delay[20]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43919), .COUT(n43920), .S0(n77[19]), .S1(n77[20]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(145[31:54])
    defparam sub_31_add_2_21.INIT0 = 16'h5555;
    defparam sub_31_add_2_21.INIT1 = 16'h5555;
    defparam sub_31_add_2_21.INJECT1_0 = "NO";
    defparam sub_31_add_2_21.INJECT1_1 = "NO";
    LUT4 i26183_4_lut_4_lut (.A(n52193), .B(n63), .C(n77[23]), .D(count_wd_delay[23]), 
         .Z(count_wd_delay_31__N_1216[23])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[19:72])
    defparam i26183_4_lut_4_lut.init = 16'h5140;
    PFUMX i40636 (.BLUT(n51738), .ALUT(n51737), .C0(\i2c_top_debug[2] ), 
          .Z(n51739));
    LUT4 i26174_4_lut_4_lut (.A(n52193), .B(n63), .C(n77[29]), .D(count_wd_delay[29]), 
         .Z(count_wd_delay_31__N_1216[29])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[19:72])
    defparam i26174_4_lut_4_lut.init = 16'h5140;
    LUT4 led_data_out_4__I_0_860_Mux_0_i1_3_lut_4_lut (.A(delay_timer_at_init), 
         .B(n66), .C(\next_i2c_device_driver_state[0] ), .D(\next_i2c_state_4__N_1090[0] ), 
         .Z(n1)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C+(D)))+!A !(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam led_data_out_4__I_0_860_Mux_0_i1_3_lut_4_lut.init = 16'h7f70;
    LUT4 i25769_2_lut_3_lut (.A(delay_timer_at_init), .B(n66), .C(\next_i2c_device_driver_state[0] ), 
         .Z(n1_adj_1)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(169[14] 181[12])
    defparam i25769_2_lut_3_lut.init = 16'h8080;
    CCU2D sub_31_add_2_19 (.A0(count_wd_delay[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_wd_delay[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43918), .COUT(n43919), .S0(count_wd_delay_31__N_1300[17]), 
          .S1(n77[18]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(145[31:54])
    defparam sub_31_add_2_19.INIT0 = 16'h5555;
    defparam sub_31_add_2_19.INIT1 = 16'h5555;
    defparam sub_31_add_2_19.INJECT1_0 = "NO";
    defparam sub_31_add_2_19.INJECT1_1 = "NO";
    CCU2D sub_31_add_2_17 (.A0(count_wd_delay[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_wd_delay[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43917), .COUT(n43918), .S0(count_wd_delay_31__N_1300[15]), 
          .S1(n77[16]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(145[31:54])
    defparam sub_31_add_2_17.INIT0 = 16'h5555;
    defparam sub_31_add_2_17.INIT1 = 16'h5555;
    defparam sub_31_add_2_17.INJECT1_0 = "NO";
    defparam sub_31_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_31_add_2_15 (.A0(count_wd_delay[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_wd_delay[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43916), .COUT(n43917), .S0(n77[13]), .S1(count_wd_delay_31__N_1300[14]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(145[31:54])
    defparam sub_31_add_2_15.INIT0 = 16'h5555;
    defparam sub_31_add_2_15.INIT1 = 16'h5555;
    defparam sub_31_add_2_15.INJECT1_0 = "NO";
    defparam sub_31_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_31_add_2_13 (.A0(count_wd_delay[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_wd_delay[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43915), .COUT(n43916), .S0(count_wd_delay_31__N_1300[11]), 
          .S1(n77[12]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(145[31:54])
    defparam sub_31_add_2_13.INIT0 = 16'h5555;
    defparam sub_31_add_2_13.INIT1 = 16'h5555;
    defparam sub_31_add_2_13.INJECT1_0 = "NO";
    defparam sub_31_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_31_add_2_11 (.A0(count_wd_delay[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_wd_delay[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43914), .COUT(n43915), .S0(count_wd_delay_31__N_1300[9]), 
          .S1(n77[10]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(145[31:54])
    defparam sub_31_add_2_11.INIT0 = 16'h5555;
    defparam sub_31_add_2_11.INIT1 = 16'h5555;
    defparam sub_31_add_2_11.INJECT1_0 = "NO";
    defparam sub_31_add_2_11.INJECT1_1 = "NO";
    LUT4 i26184_4_lut_4_lut (.A(n52193), .B(n63), .C(n77[22]), .D(count_wd_delay[22]), 
         .Z(count_wd_delay_31__N_1216[22])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[19:72])
    defparam i26184_4_lut_4_lut.init = 16'h5140;
    CCU2D sub_31_add_2_9 (.A0(count_wd_delay[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_wd_delay[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43913), .COUT(n43914), .S0(n77[7]), .S1(n77[8]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(145[31:54])
    defparam sub_31_add_2_9.INIT0 = 16'h5555;
    defparam sub_31_add_2_9.INIT1 = 16'h5555;
    defparam sub_31_add_2_9.INJECT1_0 = "NO";
    defparam sub_31_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_31_add_2_7 (.A0(count_wd_delay[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_wd_delay[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43912), .COUT(n43913), .S0(n77[5]), .S1(count_wd_delay_31__N_1300[6]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(145[31:54])
    defparam sub_31_add_2_7.INIT0 = 16'h5555;
    defparam sub_31_add_2_7.INIT1 = 16'h5555;
    defparam sub_31_add_2_7.INJECT1_0 = "NO";
    defparam sub_31_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_31_add_2_5 (.A0(count_wd_delay[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_wd_delay[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43911), .COUT(n43912), .S0(n77[3]), .S1(n77[4]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(145[31:54])
    defparam sub_31_add_2_5.INIT0 = 16'h5555;
    defparam sub_31_add_2_5.INIT1 = 16'h5555;
    defparam sub_31_add_2_5.INJECT1_0 = "NO";
    defparam sub_31_add_2_5.INJECT1_1 = "NO";
    LUT4 i26185_4_lut_4_lut (.A(n52193), .B(n63), .C(n77[20]), .D(count_wd_delay[20]), 
         .Z(count_wd_delay_31__N_1216[20])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[19:72])
    defparam i26185_4_lut_4_lut.init = 16'h5140;
    LUT4 i27031_4_lut (.A(n38161), .B(\i2c_top_debug[3] ), .C(n52424), 
         .D(n53886), .Z(n15)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B+!(C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i27031_4_lut.init = 16'hcfdd;
    CCU2D sub_31_add_2_3 (.A0(count_wd_delay[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count_wd_delay[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43910), .COUT(n43911), .S0(n77[1]), .S1(n77[2]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(145[31:54])
    defparam sub_31_add_2_3.INIT0 = 16'h5555;
    defparam sub_31_add_2_3.INIT1 = 16'h5555;
    defparam sub_31_add_2_3.INJECT1_0 = "NO";
    defparam sub_31_add_2_3.INJECT1_1 = "NO";
    LUT4 i2_2_lut_rep_516 (.A(n53886), .B(\i2c_top_debug[3] ), .Z(n52452)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i2_2_lut_rep_516.init = 16'heeee;
    LUT4 i39865_2_lut_3_lut (.A(n53886), .B(\i2c_top_debug[3] ), .C(\i2c_top_debug[4] ), 
         .Z(n27058)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i39865_2_lut_3_lut.init = 16'h0101;
    CCU2D sub_31_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count_wd_delay[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n43910), .S1(n77[0]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(145[31:54])
    defparam sub_31_add_2_1.INIT0 = 16'hF000;
    defparam sub_31_add_2_1.INIT1 = 16'h5555;
    defparam sub_31_add_2_1.INJECT1_0 = "NO";
    defparam sub_31_add_2_1.INJECT1_1 = "NO";
    PFUMX i41283 (.BLUT(n53178), .ALUT(n53173), .C0(\i2c_top_debug[4] ), 
          .Z(next_i2c_cmd_state_5__N_1479[1]));
    PFUMX i41281 (.BLUT(n53176), .ALUT(n53175), .C0(\i2c_top_debug[5] ), 
          .Z(n53177));
    LUT4 i1_2_lut_rep_519 (.A(byte_wr_left[1]), .B(byte_wr_left[0]), .Z(n52455)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(750[46:65])
    defparam i1_2_lut_rep_519.init = 16'hdddd;
    LUT4 i1_2_lut_rep_292_2_lut_3_lut_4_lut (.A(byte_wr_left[1]), .B(byte_wr_left[0]), 
         .C(ack_flag), .D(ack), .Z(n52228)) /* synthesis lut_function=(!(A ((C (D))+!B)+!A (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(750[46:65])
    defparam i1_2_lut_rep_292_2_lut_3_lut_4_lut.init = 16'h0ddd;
    LUT4 i11_3_lut_4_lut (.A(byte_wr_left[1]), .B(byte_wr_left[0]), .C(\data_reg[0] ), 
         .D(\data_reg[8] ), .Z(n1296[0])) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(750[46:65])
    defparam i11_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i1_2_lut_3_lut_adj_311 (.A(byte_wr_left[1]), .B(byte_wr_left[0]), 
         .C(\data_reg[7] ), .Z(n7_adj_5239)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(750[46:65])
    defparam i1_2_lut_3_lut_adj_311.init = 16'hd0d0;
    LUT4 i26186_4_lut_4_lut (.A(n52193), .B(n63), .C(n77[19]), .D(count_wd_delay[19]), 
         .Z(count_wd_delay_31__N_1216[19])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[19:72])
    defparam i26186_4_lut_4_lut.init = 16'h5140;
    LUT4 i39825_4_lut (.A(wd_event_active), .B(n76), .C(n8_adj_5256), 
         .D(n44475), .Z(sys_clk_enable_148)) /* synthesis lut_function=(A+!(B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(267[14] 1038[12])
    defparam i39825_4_lut.init = 16'haaab;
    LUT4 i3_4_lut (.A(n49_adj_5220), .B(\i2c_top_debug[5] ), .C(n52299), 
         .D(n52436), .Z(n8_adj_5256)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(267[14] 1038[12])
    defparam i3_4_lut.init = 16'hfeee;
    LUT4 i7683_2_lut_rep_239_3_lut_4_lut (.A(byte_rd_left[3]), .B(n52239), 
         .C(byte_rd_left[5]), .D(byte_rd_left[4]), .Z(n52175)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(226[29:50])
    defparam i7683_2_lut_rep_239_3_lut_4_lut.init = 16'hfffe;
    FD1P3AX byte_wr_left_6626__i1 (.D(n17[1]), .SP(sys_clk_enable_148), 
            .CK(sys_clk), .Q(byte_wr_left[1]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(750[46:65])
    defparam byte_wr_left_6626__i1.GSR = "ENABLED";
    LUT4 i2_2_lut_rep_528 (.A(\i2c_top_debug[3] ), .B(\i2c_top_debug[4] ), 
         .Z(n52464)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i2_2_lut_rep_528.init = 16'heeee;
    PFUMX i38643 (.BLUT(n10_adj_5219), .ALUT(n14_adj_5253), .C0(n52416), 
          .Z(n49438));
    LUT4 i1_2_lut_rep_352_3_lut (.A(\i2c_top_debug[3] ), .B(\i2c_top_debug[4] ), 
         .C(\i2c_top_debug[5] ), .Z(n52288)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i1_2_lut_rep_352_3_lut.init = 16'hfefe;
    LUT4 clear_waiting_us_N_1211_I_0_2_lut (.A(clear_waiting_us), .B(resetn), 
         .Z(count_us_11__N_1215)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_device_driver.v(140[16] 159[6])
    defparam clear_waiting_us_N_1211_I_0_2_lut.init = 16'h4444;
    PFUMX i41278 (.BLUT(n22), .ALUT(n53171), .C0(\i2c_top_debug[3] ), 
          .Z(n53172));
    LUT4 i3_4_lut_adj_312 (.A(n52425), .B(n52316), .C(n52306), .D(n52318), 
         .Z(clear_waiting_us)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(254[14] 1038[12])
    defparam i3_4_lut_adj_312.init = 16'hfffe;
    LUT4 i26187_4_lut_4_lut (.A(n52193), .B(n63), .C(n77[18]), .D(count_wd_delay[18]), 
         .Z(count_wd_delay_31__N_1216[18])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[19:72])
    defparam i26187_4_lut_4_lut.init = 16'h5140;
    PFUMX i40998 (.BLUT(n52606), .ALUT(n52607), .C0(\i2c_top_debug[3] ), 
          .Z(n52608));
    LUT4 i2_3_lut_rep_257_4_lut (.A(n52318), .B(n52248), .C(n52288), .D(n52289), 
         .Z(n52193)) /* synthesis lut_function=(A+!(B (C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(254[14] 1038[12])
    defparam i2_3_lut_rep_257_4_lut.init = 16'hbbbf;
    FD1S3DX byte_rd_left_i1_19954_19955_reset (.D(byte_rd_left_5__N_1248[1]), 
            .CK(data_latch), .CD(byte_rd_left_5__N_1279), .Q(n30627)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(225[14] 227[12])
    defparam byte_rd_left_i1_19954_19955_reset.GSR = "DISABLED";
    LUT4 i26190_4_lut_4_lut (.A(n52193), .B(n63), .C(n77[16]), .D(count_wd_delay[16]), 
         .Z(count_wd_delay_31__N_1216[16])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[19:72])
    defparam i26190_4_lut_4_lut.init = 16'h5140;
    LUT4 byte_wr_left_6626_mux_6_i1_4_lut (.A(is_2_byte_reg), .B(byte_wr_left[0]), 
         .C(n6849), .D(n48107), .Z(n17[0])) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(750[46:65])
    defparam byte_wr_left_6626_mux_6_i1_4_lut.init = 16'h3530;
    LUT4 i3_4_lut_adj_313 (.A(n52140), .B(n52425), .C(n53886), .D(n37653), 
         .Z(n6849)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[14] 151[12])
    defparam i3_4_lut_adj_313.init = 16'h0080;
    LUT4 n51536_bdd_4_lut_41634 (.A(n51536), .B(n52425), .C(\i2c_top_debug[0] ), 
         .D(\i2c_top_debug[1] ), .Z(n53176)) /* synthesis lut_function=(A+!(((D)+!C)+!B)) */ ;
    defparam n51536_bdd_4_lut_41634.init = 16'haaea;
    LUT4 i1_2_lut_rep_523 (.A(byte_wr_left[1]), .B(byte_wr_left[0]), .Z(n52459)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(750[46:65])
    defparam i1_2_lut_rep_523.init = 16'heeee;
    PFUMX mux_464_Mux_2_i31 (.BLUT(n25), .ALUT(n28215), .C0(n49652), .Z(n31_adj_5248)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;
    LUT4 i1_2_lut_3_lut_4_lut_adj_314 (.A(byte_rd_left[3]), .B(n52239), 
         .C(byte_rd_left[5]), .D(byte_rd_left[4]), .Z(byte_rd_left_5__N_1248[5])) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)+!C !(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(226[29:50])
    defparam i1_2_lut_3_lut_4_lut_adj_314.init = 16'hf0e1;
    PFUMX mux_464_Mux_5_i63 (.BLUT(n48814), .ALUT(n62_adj_5221), .C0(\i2c_top_debug[5] ), 
          .Z(next_i2c_cmd_state_5__N_1479[5])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;
    L6MUX21 i38609 (.D0(n49402), .D1(n49403), .SD(\next_i2c_device_driver_state[2] ), 
            .Z(\next_data_reg_15__N_362[0] ));
    LUT4 i1_3_lut_4_lut_adj_315 (.A(byte_wr_left[1]), .B(byte_wr_left[0]), 
         .C(n53), .D(\i2c_top_debug[1] ), .Z(n50)) /* synthesis lut_function=(A (C+(D))+!A (B (C+(D))+!B (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(750[46:65])
    defparam i1_3_lut_4_lut_adj_315.init = 16'hffe0;
    PFUMX i38595 (.BLUT(n10_c), .ALUT(n14_adj_5251), .C0(n52416), .Z(n49390));
    LUT4 i3_3_lut_rep_370_4_lut (.A(\i2c_top_debug[3] ), .B(\i2c_top_debug[4] ), 
         .C(n53886), .D(\i2c_top_debug[5] ), .Z(n52306)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(268[13] 1037[20])
    defparam i3_3_lut_rep_370_4_lut.init = 16'hfffe;
    LUT4 i26193_4_lut_4_lut (.A(n52193), .B(n63), .C(n77[10]), .D(count_wd_delay[10]), 
         .Z(count_wd_delay_31__N_1216[10])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[19:72])
    defparam i26193_4_lut_4_lut.init = 16'h5140;
    PFUMX i40952 (.BLUT(n52537), .ALUT(n52538), .C0(\i2c_top_debug[3] ), 
          .Z(n52539));
    LUT4 i2_3_lut_4_lut_adj_316 (.A(byte_wr_left[1]), .B(byte_wr_left[0]), 
         .C(\i2c_top_debug[0] ), .D(\i2c_top_debug[1] ), .Z(n48845)) /* synthesis lut_function=(A (C+(D))+!A ((C+(D))+!B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(750[46:65])
    defparam i2_3_lut_4_lut_adj_316.init = 16'hfff1;
    PFUMX i38624 (.BLUT(n49417), .ALUT(n49418), .C0(\i2c_top_debug[4] ), 
          .Z(n49419));
    PFUMX i2c_top_debug_5__I_0_767_Mux_0_i63 (.BLUT(n49767), .ALUT(n49768), 
          .C0(n49672), .Z(next_addr_7__N_1160[0])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;
    LUT4 i7029_1_lut_rep_238_3_lut_4_lut (.A(n52318), .B(n52248), .C(n52288), 
         .D(n52289), .Z(n52174)) /* synthesis lut_function=(!(A+!(B (C+(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(254[14] 1038[12])
    defparam i7029_1_lut_rep_238_3_lut_4_lut.init = 16'h4440;
    LUT4 i26191_4_lut_4_lut (.A(n52193), .B(n63), .C(n77[13]), .D(count_wd_delay[13]), 
         .Z(count_wd_delay_31__N_1216[13])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[19:72])
    defparam i26191_4_lut_4_lut.init = 16'h5140;
    FD1P3JX count_wd_delay_i6 (.D(count_wd_delay_31__N_1300[6]), .SP(sys_clk_enable_231), 
            .PD(n52193), .CK(sys_clk), .Q(count_wd_delay[6])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[14] 151[12])
    defparam count_wd_delay_i6.GSR = "ENABLED";
    FD1P3JX count_wd_delay_i9 (.D(count_wd_delay_31__N_1300[9]), .SP(sys_clk_enable_231), 
            .PD(n52193), .CK(sys_clk), .Q(count_wd_delay[9])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[14] 151[12])
    defparam count_wd_delay_i9.GSR = "ENABLED";
    FD1P3JX count_wd_delay_i11 (.D(count_wd_delay_31__N_1300[11]), .SP(sys_clk_enable_231), 
            .PD(n52193), .CK(sys_clk), .Q(count_wd_delay[11])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[14] 151[12])
    defparam count_wd_delay_i11.GSR = "ENABLED";
    FD1P3JX count_wd_delay_i14 (.D(count_wd_delay_31__N_1300[14]), .SP(sys_clk_enable_231), 
            .PD(n52193), .CK(sys_clk), .Q(count_wd_delay[14])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[14] 151[12])
    defparam count_wd_delay_i14.GSR = "ENABLED";
    FD1P3JX count_wd_delay_i15 (.D(count_wd_delay_31__N_1300[15]), .SP(sys_clk_enable_231), 
            .PD(n52193), .CK(sys_clk), .Q(count_wd_delay[15])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[14] 151[12])
    defparam count_wd_delay_i15.GSR = "ENABLED";
    FD1P3JX count_wd_delay_i17 (.D(count_wd_delay_31__N_1300[17]), .SP(sys_clk_enable_231), 
            .PD(n52193), .CK(sys_clk), .Q(count_wd_delay[17])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[14] 151[12])
    defparam count_wd_delay_i17.GSR = "ENABLED";
    FD1P3JX count_wd_delay_i21 (.D(count_wd_delay_31__N_1300[21]), .SP(sys_clk_enable_231), 
            .PD(n52193), .CK(sys_clk), .Q(count_wd_delay[21])) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(140[14] 151[12])
    defparam count_wd_delay_i21.GSR = "ENABLED";
    FD1S1I next_we_I_0 (.D(n52300), .CK(next_addr_7__N_1168), .CD(n51040), 
           .Q(next_we)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(231[5] 1039[8])
    defparam next_we_I_0.GSR = "DISABLED";
    FD1S3BX byte_rd_left_i1_19954_19955_set (.D(byte_rd_left_5__N_1248[1]), 
            .CK(data_latch), .PD(byte_rd_left_5__N_1265), .Q(n30626)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(225[14] 227[12])
    defparam byte_rd_left_i1_19954_19955_set.GSR = "DISABLED";
    FD1S3DX byte_rd_left_i0_19950_19951_reset (.D(n52439), .CK(data_latch), 
            .CD(byte_rd_left_5__N_1282), .Q(n30623)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(225[14] 227[12])
    defparam byte_rd_left_i0_19950_19951_reset.GSR = "DISABLED";
    FD1S3BX byte_rd_left_i0_19950_19951_set (.D(n52439), .CK(data_latch), 
            .PD(byte_rd_left_5__N_1266), .Q(n30622)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(225[14] 227[12])
    defparam byte_rd_left_i0_19950_19951_set.GSR = "DISABLED";
    FD1S3DX count_us_i0_i0_19938_19939_reset (.D(n26[0]), .CK(sys_clk), 
            .CD(count_us_11__N_1215), .Q(n30611)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(128[14] 131[34])
    defparam count_us_i0_i0_19938_19939_reset.GSR = "DISABLED";
    FD1S3DX count_us_i0_i6_19935_19936_reset (.D(n26[6]), .CK(sys_clk), 
            .CD(count_us_11__N_1215), .Q(n30608)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(128[14] 131[34])
    defparam count_us_i0_i6_19935_19936_reset.GSR = "DISABLED";
    FD1S3DX count_us_i0_i8_19932_19933_reset (.D(n26[8]), .CK(sys_clk), 
            .CD(count_us_11__N_1215), .Q(n30605)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(128[14] 131[34])
    defparam count_us_i0_i8_19932_19933_reset.GSR = "DISABLED";
    FD1S3DX count_us_i0_i9_19929_19930_reset (.D(n26[9]), .CK(sys_clk), 
            .CD(count_us_11__N_1215), .Q(n30602)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(128[14] 131[34])
    defparam count_us_i0_i9_19929_19930_reset.GSR = "DISABLED";
    FD1S3DX count_us_i0_i10_19926_19927_reset (.D(n26[10]), .CK(sys_clk), 
            .CD(count_us_11__N_1215), .Q(n30599)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(128[14] 131[34])
    defparam count_us_i0_i10_19926_19927_reset.GSR = "DISABLED";
    FD1S3DX count_us_i0_i11_19923_19924_reset (.D(n26[11]), .CK(sys_clk), 
            .CD(count_us_11__N_1215), .Q(n30596)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(128[14] 131[34])
    defparam count_us_i0_i11_19923_19924_reset.GSR = "DISABLED";
    FD1S3AY count_us_i0_i11_19923_19924_set (.D(n26[11]), .CK(sys_clk), 
            .Q(n30595)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(128[14] 131[34])
    defparam count_us_i0_i11_19923_19924_set.GSR = "ENABLED";
    PFUMX i2c_top_debug_5__I_0_768_Mux_0_i31 (.BLUT(n48098), .ALUT(n30), 
          .C0(\i2c_top_debug[4] ), .Z(n31)) /* synthesis LSE_LINE_FILE_ID=30, LSE_LCOL=16, LSE_RCOL=6, LSE_LLINE=140, LSE_RLINE=159 */ ;
    I2C_EFB_WB data_rx_7__I_0 (.sys_clk(sys_clk), .data_rx_7__N_1159(data_rx_7__N_1159), 
            .stb(stb), .we(we), .GND_net(GND_net), .\addr[2] (addr[2]), 
            .\addr[1] (addr[1]), .\addr[0] (addr[0]), .data_tx({data_tx_c}), 
            .data_rx({data_rx_adj_5257}), .ack(ack), .i2c2_sdaoen(i2c2_sdaoen), 
            .i2c2_sdao(i2c2_sdao), .i2c2_scloen(i2c2_scloen), .i2c2_sclo(i2c2_sclo), 
            .i2c2_sdai(i2c2_sdai), .i2c2_scli(i2c2_scli), .i2c1_sdaoen(i2c1_sdaoen), 
            .i2c1_sdao(i2c1_sdao), .i2c1_scloen(i2c1_scloen), .i2c1_sclo(i2c1_sclo), 
            .i2c1_sdai(i2c1_sdai), .i2c1_scli(i2c1_scli), .VCC_net(VCC_net), 
            .n53(n53), .n52466(n52466), .ack_flag(ack_flag), .n52301(n52301)) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(99[16] 115[2])
    
endmodule
//
// Verilog Description of module I2C_EFB_WB
//

module I2C_EFB_WB (sys_clk, data_rx_7__N_1159, stb, we, GND_net, \addr[2] , 
            \addr[1] , \addr[0] , data_tx, data_rx, ack, i2c2_sdaoen, 
            i2c2_sdao, i2c2_scloen, i2c2_sclo, i2c2_sdai, i2c2_scli, 
            i2c1_sdaoen, i2c1_sdao, i2c1_scloen, i2c1_sclo, i2c1_sdai, 
            i2c1_scli, VCC_net, n53, n52466, ack_flag, n52301) /* synthesis NGD_DRC_MASK=1, syn_module_defined=1 */ ;
    input sys_clk;
    input data_rx_7__N_1159;
    input stb;
    input we;
    input GND_net;
    input \addr[2] ;
    input \addr[1] ;
    input \addr[0] ;
    input [7:0]data_tx;
    output [7:0]data_rx;
    output ack;
    output i2c2_sdaoen;
    output i2c2_sdao;
    output i2c2_scloen;
    output i2c2_sclo;
    input i2c2_sdai;
    input i2c2_scli;
    output i2c1_sdaoen;
    output i2c1_sdao;
    output i2c1_scloen;
    output i2c1_sclo;
    input i2c1_sdai;
    input i2c1_scli;
    input VCC_net;
    output n53;
    output n52466;
    input ack_flag;
    output n52301;
    
    wire sys_clk /* synthesis SET_AS_NETWORK=sys_clk, is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(220[10:17])
    wire i2c2_scli /* synthesis is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_efb_wb.v(34[10:19])
    wire i2c1_scli /* synthesis is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_efb_wb.v(40[10:19])
    
    EFB EFBInst_0 (.WBCLKI(sys_clk), .WBRSTI(data_rx_7__N_1159), .WBCYCI(stb), 
        .WBSTBI(stb), .WBWEI(we), .WBADRI0(\addr[0] ), .WBADRI1(\addr[1] ), 
        .WBADRI2(\addr[2] ), .WBADRI3(GND_net), .WBADRI4(GND_net), .WBADRI5(GND_net), 
        .WBADRI6(stb), .WBADRI7(GND_net), .WBDATI0(data_tx[0]), .WBDATI1(data_tx[1]), 
        .WBDATI2(data_tx[2]), .WBDATI3(data_tx[3]), .WBDATI4(data_tx[4]), 
        .WBDATI5(data_tx[5]), .WBDATI6(data_tx[6]), .WBDATI7(data_tx[7]), 
        .I2C1SCLI(i2c1_scli), .I2C1SDAI(i2c1_sdai), .I2C2SCLI(i2c2_scli), 
        .I2C2SDAI(i2c2_sdai), .SPISCKI(GND_net), .SPIMISOI(GND_net), .SPIMOSII(GND_net), 
        .SPISCSN(GND_net), .TCCLKI(GND_net), .TCRSTN(GND_net), .TCIC(GND_net), 
        .UFMSN(VCC_net), .PLL0DATI0(GND_net), .PLL0DATI1(GND_net), .PLL0DATI2(GND_net), 
        .PLL0DATI3(GND_net), .PLL0DATI4(GND_net), .PLL0DATI5(GND_net), 
        .PLL0DATI6(GND_net), .PLL0DATI7(GND_net), .PLL0ACKI(GND_net), 
        .PLL1DATI0(GND_net), .PLL1DATI1(GND_net), .PLL1DATI2(GND_net), 
        .PLL1DATI3(GND_net), .PLL1DATI4(GND_net), .PLL1DATI5(GND_net), 
        .PLL1DATI6(GND_net), .PLL1DATI7(GND_net), .PLL1ACKI(GND_net), 
        .WBDATO0(data_rx[0]), .WBDATO1(data_rx[1]), .WBDATO2(data_rx[2]), 
        .WBDATO3(data_rx[3]), .WBDATO4(data_rx[4]), .WBDATO5(data_rx[5]), 
        .WBDATO6(data_rx[6]), .WBDATO7(data_rx[7]), .WBACKO(ack), .I2C1SCLO(i2c1_sclo), 
        .I2C1SCLOEN(i2c1_scloen), .I2C1SDAO(i2c1_sdao), .I2C1SDAOEN(i2c1_sdaoen), 
        .I2C2SCLO(i2c2_sclo), .I2C2SCLOEN(i2c2_scloen), .I2C2SDAO(i2c2_sdao), 
        .I2C2SDAOEN(i2c2_sdaoen)) /* synthesis syn_instantiated=1, LSE_LINE_FILE_ID=8, LSE_LCOL=16, LSE_RCOL=2, LSE_LLINE=99, LSE_RLINE=115 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(99[16] 115[2])
    defparam EFBInst_0.EFB_I2C1 = "ENABLED";
    defparam EFBInst_0.EFB_I2C2 = "ENABLED";
    defparam EFBInst_0.EFB_SPI = "DISABLED";
    defparam EFBInst_0.EFB_TC = "DISABLED";
    defparam EFBInst_0.EFB_TC_PORTMODE = "WB";
    defparam EFBInst_0.EFB_UFM = "DISABLED";
    defparam EFBInst_0.EFB_WB_CLK_FREQ = "38.0";
    defparam EFBInst_0.DEV_DENSITY = "6900L";
    defparam EFBInst_0.UFM_INIT_PAGES = 0;
    defparam EFBInst_0.UFM_INIT_START_PAGE = 0;
    defparam EFBInst_0.UFM_INIT_ALL_ZEROS = "ENABLED";
    defparam EFBInst_0.UFM_INIT_FILE_NAME = "NONE";
    defparam EFBInst_0.UFM_INIT_FILE_FORMAT = "HEX";
    defparam EFBInst_0.I2C1_ADDRESSING = "7BIT";
    defparam EFBInst_0.I2C2_ADDRESSING = "7BIT";
    defparam EFBInst_0.I2C1_SLAVE_ADDR = "0b1000001";
    defparam EFBInst_0.I2C2_SLAVE_ADDR = "0b1000010";
    defparam EFBInst_0.I2C1_BUS_PERF = "400kHz";
    defparam EFBInst_0.I2C2_BUS_PERF = "400kHz";
    defparam EFBInst_0.I2C1_CLK_DIVIDER = 24;
    defparam EFBInst_0.I2C2_CLK_DIVIDER = 24;
    defparam EFBInst_0.I2C1_GEN_CALL = "DISABLED";
    defparam EFBInst_0.I2C2_GEN_CALL = "DISABLED";
    defparam EFBInst_0.I2C1_WAKEUP = "DISABLED";
    defparam EFBInst_0.I2C2_WAKEUP = "DISABLED";
    defparam EFBInst_0.SPI_MODE = "MASTER";
    defparam EFBInst_0.SPI_CLK_DIVIDER = 1;
    defparam EFBInst_0.SPI_LSB_FIRST = "DISABLED";
    defparam EFBInst_0.SPI_CLK_INV = "DISABLED";
    defparam EFBInst_0.SPI_PHASE_ADJ = "DISABLED";
    defparam EFBInst_0.SPI_SLAVE_HANDSHAKE = "DISABLED";
    defparam EFBInst_0.SPI_INTR_TXRDY = "DISABLED";
    defparam EFBInst_0.SPI_INTR_RXRDY = "DISABLED";
    defparam EFBInst_0.SPI_INTR_TXOVR = "DISABLED";
    defparam EFBInst_0.SPI_INTR_RXOVR = "DISABLED";
    defparam EFBInst_0.SPI_WAKEUP = "DISABLED";
    defparam EFBInst_0.TC_MODE = "CTCM";
    defparam EFBInst_0.TC_SCLK_SEL = "PCLOCK";
    defparam EFBInst_0.TC_CCLK_SEL = 1;
    defparam EFBInst_0.GSR = "ENABLED";
    defparam EFBInst_0.TC_TOP_SET = 65535;
    defparam EFBInst_0.TC_OCR_SET = 32767;
    defparam EFBInst_0.TC_OC_MODE = "TOGGLE";
    defparam EFBInst_0.TC_RESETN = "ENABLED";
    defparam EFBInst_0.TC_TOP_SEL = "OFF";
    defparam EFBInst_0.TC_OV_INT = "OFF";
    defparam EFBInst_0.TC_OCR_INT = "OFF";
    defparam EFBInst_0.TC_ICR_INT = "OFF";
    defparam EFBInst_0.TC_OVERFLOW = "DISABLED";
    defparam EFBInst_0.TC_ICAPTURE = "DISABLED";
    LUT4 i1_2_lut (.A(data_rx[6]), .B(data_rx[2]), .Z(n53)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(99[16] 115[2])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i1_2_lut_rep_530 (.A(data_rx[2]), .B(data_rx[5]), .Z(n52466)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(99[16] 115[2])
    defparam i1_2_lut_rep_530.init = 16'hdddd;
    LUT4 i1_2_lut_rep_365_3_lut_4_lut (.A(data_rx[2]), .B(data_rx[5]), .C(ack_flag), 
         .D(ack), .Z(n52301)) /* synthesis lut_function=((B+!(C (D)))+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/i2c_module_top.v(99[16] 115[2])
    defparam i1_2_lut_rep_365_3_lut_4_lut.init = 16'hdfff;
    
endmodule
//
// Verilog Description of module z_linear_velocity_comp
//

module z_linear_velocity_comp (n53884, sys_clk, \next_state_4__N_1567[2] , 
            \z_linear_velocity[3] , \z_linear_velocity[1] , \z_linear_velocity[2] , 
            n50715, \z_linear_velocity[6] , \z_linear_velocity[5] , \z_linear_velocity[7] , 
            \z_linear_velocity[4] , n43332, GND_net, \tx_byte_index[0] , 
            \tx_byte_index[1] , n52168, n43302, n43303, n27734, n48081, 
            n123, n52255, \next_dat_i_15__N_4452[3] , \next_state_4__N_1656[2] , 
            us_clk_enable_103, n46653, n52341, n37731, n52342, n15182, 
            \state[2] , \state[5] , n43309, \z_linear_velocity[10] , 
            \z_linear_velocity[11] , \VL53L1X_range_mm[1] , \VL53L1X_range_mm[2] , 
            \VL53L1X_range_mm[3] , \VL53L1X_range_mm[4] , \VL53L1X_range_mm[5] , 
            \VL53L1X_range_mm[6] , \VL53L1X_range_mm[7] , \VL53L1X_range_mm[8] , 
            \VL53L1X_range_mm[9] , \VL53L1X_range_mm[10] , \VL53L1X_range_mm[11] , 
            \VL53L1X_range_mm[12] , \VL53L1X_range_mm[13] , \VL53L1X_range_mm[14] , 
            \z_linear_velocity[12] , \z_linear_velocity[13] , \z_linear_velocity[14] , 
            \z_linear_velocity[15] , \VL53L1X_range_mm[0] , \z_linear_velocity[8] , 
            \z_linear_velocity[9] ) /* synthesis syn_module_defined=1 */ ;
    input n53884;
    input sys_clk;
    input \next_state_4__N_1567[2] ;
    output \z_linear_velocity[3] ;
    output \z_linear_velocity[1] ;
    output \z_linear_velocity[2] ;
    output n50715;
    output \z_linear_velocity[6] ;
    output \z_linear_velocity[5] ;
    output \z_linear_velocity[7] ;
    output \z_linear_velocity[4] ;
    output n43332;
    input GND_net;
    input \tx_byte_index[0] ;
    input \tx_byte_index[1] ;
    output n52168;
    output n43302;
    output n43303;
    input n27734;
    input n48081;
    input n123;
    input n52255;
    output \next_dat_i_15__N_4452[3] ;
    input \next_state_4__N_1656[2] ;
    input us_clk_enable_103;
    output n46653;
    input n52341;
    input n37731;
    input n52342;
    output n15182;
    input \state[2] ;
    input \state[5] ;
    output n43309;
    output \z_linear_velocity[10] ;
    output \z_linear_velocity[11] ;
    input \VL53L1X_range_mm[1] ;
    input \VL53L1X_range_mm[2] ;
    input \VL53L1X_range_mm[3] ;
    input \VL53L1X_range_mm[4] ;
    input \VL53L1X_range_mm[5] ;
    input \VL53L1X_range_mm[6] ;
    input \VL53L1X_range_mm[7] ;
    input \VL53L1X_range_mm[8] ;
    input \VL53L1X_range_mm[9] ;
    input \VL53L1X_range_mm[10] ;
    input \VL53L1X_range_mm[11] ;
    input \VL53L1X_range_mm[12] ;
    input \VL53L1X_range_mm[13] ;
    input \VL53L1X_range_mm[14] ;
    output \z_linear_velocity[12] ;
    output \z_linear_velocity[13] ;
    output \z_linear_velocity[14] ;
    output \z_linear_velocity[15] ;
    input \VL53L1X_range_mm[0] ;
    output \z_linear_velocity[8] ;
    output \z_linear_velocity[9] ;
    
    wire next_state_4__N_1576 /* synthesis is_clock=1, SET_AS_NETWORK=\ZLV/next_state_4__N_1576 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(48[38:48])
    wire sys_clk /* synthesis SET_AS_NETWORK=sys_clk, is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(220[10:17])
    wire [4:0]next_state;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(48[38:48])
    wire [4:0]state;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(48[31:36])
    
    wire next_state_4__N_1572, start_signal_N_1872, n49081, n52238, 
        next_state_4__N_1564, n52490, n52489, n52433, n17, n48369, 
        n50468, n48192, n52387, n43864;
    wire [10:0]n21358;
    wire [15:0]n117;
    wire [22:0]next_z_linear_velocity_calc_15__N_1577;
    
    wire n43863, n43862, n43861, n51189, n51188, n43860, n43858, 
        n8, sys_clk_enable_257, n30639, n43857, sys_clk_enable_252, 
        n27, sys_clk_enable_251, n30732, n43856, n43855, n43854, 
        n52285, n30748, n22, n43841;
    wire [15:0]z_altitude_mm_previous;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(43[37:59])
    wire [15:0]z_altitude_mm_latched;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(41[37:58])
    
    wire n43840, n43839, n43838, n43837, n43836, n43835;
    
    FD1S1AY next_state_4__I_0_i1 (.D(n53884), .CK(next_state_4__N_1576), 
            .Q(next_state[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(67[5] 82[8])
    defparam next_state_4__I_0_i1.GSR = "ENABLED";
    FD1S3AY state_i0 (.D(next_state[0]), .CK(sys_clk), .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam state_i0.GSR = "ENABLED";
    FD1S1A next_state_4__I_0_i2 (.D(next_state_4__N_1572), .CK(next_state_4__N_1576), 
           .Q(next_state[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(67[5] 82[8])
    defparam next_state_4__I_0_i2.GSR = "ENABLED";
    FD1S1I next_state_4__I_0_i3 (.D(n49081), .CK(next_state_4__N_1576), 
           .CD(start_signal_N_1872), .Q(next_state[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(67[5] 82[8])
    defparam next_state_4__I_0_i3.GSR = "ENABLED";
    FD1S1A next_state_4__I_0_i4 (.D(n52238), .CK(next_state_4__N_1576), 
           .Q(next_state[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(67[5] 82[8])
    defparam next_state_4__I_0_i4.GSR = "ENABLED";
    FD1S1A next_state_4__I_0_i5 (.D(next_state_4__N_1564), .CK(next_state_4__N_1576), 
           .Q(next_state[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(67[5] 82[8])
    defparam next_state_4__I_0_i5.GSR = "ENABLED";
    LUT4 i1_4_lut_then_3_lut_4_lut (.A(state[0]), .B(state[4]), .C(state[3]), 
         .D(state[1]), .Z(n52490)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i1_4_lut_then_3_lut_4_lut.init = 16'h0001;
    LUT4 i1_4_lut_else_3_lut_4_lut (.A(state[4]), .B(state[0]), .C(state[1]), 
         .D(state[3]), .Z(n52489)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (B (C+(D))+!B (C (D)+!C !(D))))) */ ;
    defparam i1_4_lut_else_3_lut_4_lut.init = 16'h0116;
    LUT4 i39661_3_lut_rep_302_4_lut (.A(state[0]), .B(n52433), .C(state[1]), 
         .D(state[2]), .Z(n52238)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam i39661_3_lut_rep_302_4_lut.init = 16'h0100;
    LUT4 i2_3_lut_4_lut (.A(state[0]), .B(n52433), .C(state[2]), .D(state[1]), 
         .Z(n49081)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam i2_3_lut_4_lut.init = 16'h0100;
    LUT4 i1_4_lut (.A(n17), .B(n48369), .C(n50468), .D(state[4]), .Z(next_state_4__N_1572)) /* synthesis lut_function=(!(A (B+(C (D)))+!A (B+(C+!(D))))) */ ;
    defparam i1_4_lut.init = 16'h0322;
    LUT4 i34_3_lut (.A(state[0]), .B(\next_state_4__N_1567[2] ), .C(state[1]), 
         .Z(n17)) /* synthesis lut_function=(!(A (C)+!A (B+!(C)))) */ ;
    defparam i34_3_lut.init = 16'h1a1a;
    LUT4 i37585_2_lut (.A(state[3]), .B(state[2]), .Z(n48369)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i37585_2_lut.init = 16'heeee;
    LUT4 i1_rep_74_2_lut (.A(state[1]), .B(state[0]), .Z(n50468)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_rep_74_2_lut.init = 16'heeee;
    LUT4 start_signal_I_0_448_1_lut (.A(\next_state_4__N_1567[2] ), .Z(start_signal_N_1872)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(100[17:30])
    defparam start_signal_I_0_448_1_lut.init = 16'h5555;
    LUT4 z_linear_velocity_3__bdd_3_lut_39999 (.A(\z_linear_velocity[3] ), 
         .B(\z_linear_velocity[1] ), .C(\z_linear_velocity[2] ), .Z(n50715)) /* synthesis lut_function=(A (B (C))+!A (C)) */ ;
    defparam z_linear_velocity_3__bdd_3_lut_39999.init = 16'hd0d0;
    LUT4 i39756_3_lut (.A(state[4]), .B(n48192), .C(state[3]), .Z(next_state_4__N_1564)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(107[17:27])
    defparam i39756_3_lut.init = 16'h1010;
    LUT4 i2_3_lut (.A(state[2]), .B(state[1]), .C(state[0]), .Z(n48192)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_rep_451 (.A(\z_linear_velocity[6] ), .B(\z_linear_velocity[5] ), 
         .Z(n52387)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(234[17:34])
    defparam i1_2_lut_rep_451.init = 16'heeee;
    LUT4 i14_3_lut_4_lut (.A(\z_linear_velocity[6] ), .B(\z_linear_velocity[5] ), 
         .C(\z_linear_velocity[7] ), .D(\z_linear_velocity[4] ), .Z(n43332)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B !(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(234[17:34])
    defparam i14_3_lut_4_lut.init = 16'h1fe0;
    CCU2D add_11137_12 (.A0(n21358[9]), .B0(n117[13]), .C0(GND_net), .D0(GND_net), 
          .A1(n21358[10]), .B1(n117[14]), .C1(GND_net), .D1(GND_net), 
          .CIN(n43864), .S0(next_z_linear_velocity_calc_15__N_1577[14]), 
          .S1(next_z_linear_velocity_calc_15__N_1577[15]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(108[51:107])
    defparam add_11137_12.INIT0 = 16'h5666;
    defparam add_11137_12.INIT1 = 16'h5666;
    defparam add_11137_12.INJECT1_0 = "NO";
    defparam add_11137_12.INJECT1_1 = "NO";
    CCU2D add_11137_10 (.A0(n21358[7]), .B0(n117[11]), .C0(GND_net), .D0(GND_net), 
          .A1(n21358[8]), .B1(n117[12]), .C1(GND_net), .D1(GND_net), 
          .CIN(n43863), .COUT(n43864), .S0(next_z_linear_velocity_calc_15__N_1577[12]), 
          .S1(next_z_linear_velocity_calc_15__N_1577[13]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(108[51:107])
    defparam add_11137_10.INIT0 = 16'h5666;
    defparam add_11137_10.INIT1 = 16'h5666;
    defparam add_11137_10.INJECT1_0 = "NO";
    defparam add_11137_10.INJECT1_1 = "NO";
    CCU2D add_11137_8 (.A0(n21358[5]), .B0(n117[9]), .C0(GND_net), .D0(GND_net), 
          .A1(n21358[6]), .B1(n117[10]), .C1(GND_net), .D1(GND_net), 
          .CIN(n43862), .COUT(n43863), .S0(next_z_linear_velocity_calc_15__N_1577[10]), 
          .S1(next_z_linear_velocity_calc_15__N_1577[11]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(108[51:107])
    defparam add_11137_8.INIT0 = 16'h5666;
    defparam add_11137_8.INIT1 = 16'h5666;
    defparam add_11137_8.INJECT1_0 = "NO";
    defparam add_11137_8.INJECT1_1 = "NO";
    FD1S3AX state_i4 (.D(next_state[4]), .CK(sys_clk), .Q(state[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam state_i4.GSR = "ENABLED";
    FD1S3AX state_i3 (.D(next_state[3]), .CK(sys_clk), .Q(state[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam state_i3.GSR = "ENABLED";
    FD1S3AX state_i2 (.D(next_state[2]), .CK(sys_clk), .Q(state[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam state_i2.GSR = "ENABLED";
    FD1S3AX state_i1 (.D(next_state[1]), .CK(sys_clk), .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam state_i1.GSR = "ENABLED";
    CCU2D add_11137_6 (.A0(n21358[3]), .B0(n117[7]), .C0(GND_net), .D0(GND_net), 
          .A1(n21358[4]), .B1(n117[8]), .C1(GND_net), .D1(GND_net), 
          .CIN(n43861), .COUT(n43862), .S0(next_z_linear_velocity_calc_15__N_1577[8]), 
          .S1(next_z_linear_velocity_calc_15__N_1577[9]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(108[51:107])
    defparam add_11137_6.INIT0 = 16'h5666;
    defparam add_11137_6.INIT1 = 16'h5666;
    defparam add_11137_6.INJECT1_0 = "NO";
    defparam add_11137_6.INJECT1_1 = "NO";
    LUT4 n51189_bdd_4_lut (.A(n51189), .B(n51188), .C(\tx_byte_index[0] ), 
         .D(\tx_byte_index[1] ), .Z(n52168)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C+(D))+!B (D))) */ ;
    defparam n51189_bdd_4_lut.init = 16'hffca;
    CCU2D add_11137_4 (.A0(n21358[1]), .B0(n117[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n21358[2]), .B1(n117[6]), .C1(GND_net), .D1(GND_net), 
          .CIN(n43860), .COUT(n43861), .S0(next_z_linear_velocity_calc_15__N_1577[6]), 
          .S1(next_z_linear_velocity_calc_15__N_1577[7]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(108[51:107])
    defparam add_11137_4.INIT0 = 16'h5666;
    defparam add_11137_4.INIT1 = 16'h5666;
    defparam add_11137_4.INJECT1_0 = "NO";
    defparam add_11137_4.INJECT1_1 = "NO";
    LUT4 i1_3_lut (.A(\z_linear_velocity[1] ), .B(\z_linear_velocity[3] ), 
         .C(\z_linear_velocity[2] ), .Z(n43302)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(234[17:34])
    defparam i1_3_lut.init = 16'hc8c8;
    CCU2D add_11137_2 (.A0(next_z_linear_velocity_calc_15__N_1577[1]), .B0(n117[3]), 
          .C0(GND_net), .D0(GND_net), .A1(next_z_linear_velocity_calc_15__N_1577[1]), 
          .B1(next_z_linear_velocity_calc_15__N_1577[2]), .C1(n117[4]), 
          .D1(GND_net), .COUT(n43860), .S1(next_z_linear_velocity_calc_15__N_1577[5]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(108[51:107])
    defparam add_11137_2.INIT0 = 16'h7000;
    defparam add_11137_2.INIT1 = 16'h9696;
    defparam add_11137_2.INJECT1_0 = "NO";
    defparam add_11137_2.INJECT1_1 = "NO";
    CCU2D add_11128_12 (.A0(n117[10]), .B0(n117[11]), .C0(GND_net), .D0(GND_net), 
          .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), .CIN(n43858), 
          .S0(n21358[10]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(108[51:107])
    defparam add_11128_12.INIT0 = 16'h5666;
    defparam add_11128_12.INIT1 = 16'h0000;
    defparam add_11128_12.INJECT1_0 = "NO";
    defparam add_11128_12.INJECT1_1 = "NO";
    LUT4 z_linear_velocity_2__bdd_3_lut_40283 (.A(\z_linear_velocity[2] ), 
         .B(\z_linear_velocity[3] ), .C(\z_linear_velocity[1] ), .Z(n51188)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam z_linear_velocity_2__bdd_3_lut_40283.init = 16'h0404;
    LUT4 z_linear_velocity_2__bdd_3_lut (.A(\z_linear_velocity[5] ), .B(\z_linear_velocity[6] ), 
         .C(\z_linear_velocity[7] ), .Z(n51189)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam z_linear_velocity_2__bdd_3_lut.init = 16'h1010;
    LUT4 i32721_4_lut (.A(n52387), .B(n43302), .C(\tx_byte_index[0] ), 
         .D(\z_linear_velocity[7] ), .Z(n43303)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(96[17:30])
    defparam i32721_4_lut.init = 16'hcac0;
    LUT4 i2_3_lut_rep_287 (.A(state[2]), .B(n8), .C(state[1]), .Z(sys_clk_enable_257)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i2_3_lut_rep_287.init = 16'h0404;
    LUT4 i20090_2_lut_4_lut (.A(state[2]), .B(n8), .C(state[1]), .D(next_state_4__N_1564), 
         .Z(n30639)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i20090_2_lut_4_lut.init = 16'h0004;
    CCU2D add_11128_10 (.A0(n117[8]), .B0(n117[9]), .C0(GND_net), .D0(GND_net), 
          .A1(n117[9]), .B1(n117[10]), .C1(GND_net), .D1(GND_net), .CIN(n43857), 
          .COUT(n43858), .S0(n21358[8]), .S1(n21358[9]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(108[51:107])
    defparam add_11128_10.INIT0 = 16'h5666;
    defparam add_11128_10.INIT1 = 16'h5666;
    defparam add_11128_10.INJECT1_0 = "NO";
    defparam add_11128_10.INJECT1_1 = "NO";
    LUT4 i2_4_lut (.A(n52433), .B(state[2]), .C(state[1]), .D(state[0]), 
         .Z(sys_clk_enable_252)) /* synthesis lut_function=(!(A+(B (C+(D))+!B (C+!(D))))) */ ;
    defparam i2_4_lut.init = 16'h0104;
    LUT4 i3_4_lut (.A(n27), .B(state[2]), .C(state[3]), .D(state[1]), 
         .Z(sys_clk_enable_251)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i3_4_lut.init = 16'h0002;
    LUT4 i20073_4_lut (.A(sys_clk_enable_251), .B(state[3]), .C(state[4]), 
         .D(n48192), .Z(n30732)) /* synthesis lut_function=(A (B+((D)+!C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam i20073_4_lut.init = 16'haa8a;
    CCU2D add_11128_8 (.A0(n117[6]), .B0(n117[7]), .C0(GND_net), .D0(GND_net), 
          .A1(n117[7]), .B1(n117[8]), .C1(GND_net), .D1(GND_net), .CIN(n43856), 
          .COUT(n43857), .S0(n21358[6]), .S1(n21358[7]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(108[51:107])
    defparam add_11128_8.INIT0 = 16'h5666;
    defparam add_11128_8.INIT1 = 16'h5666;
    defparam add_11128_8.INJECT1_0 = "NO";
    defparam add_11128_8.INJECT1_1 = "NO";
    LUT4 i1_4_lut_adj_279 (.A(n27734), .B(n48081), .C(n123), .D(n52255), 
         .Z(\next_dat_i_15__N_4452[3] )) /* synthesis lut_function=(A (B)+!A !(((D)+!C)+!B)) */ ;
    defparam i1_4_lut_adj_279.init = 16'h88c8;
    CCU2D add_11128_6 (.A0(n117[4]), .B0(n117[5]), .C0(GND_net), .D0(GND_net), 
          .A1(n117[5]), .B1(n117[6]), .C1(GND_net), .D1(GND_net), .CIN(n43855), 
          .COUT(n43856), .S0(n21358[4]), .S1(n21358[5]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(108[51:107])
    defparam add_11128_6.INIT0 = 16'h5666;
    defparam add_11128_6.INIT1 = 16'h5666;
    defparam add_11128_6.INJECT1_0 = "NO";
    defparam add_11128_6.INJECT1_1 = "NO";
    CCU2D add_11128_4 (.A0(next_z_linear_velocity_calc_15__N_1577[3]), .B0(n117[3]), 
          .C0(GND_net), .D0(GND_net), .A1(n117[3]), .B1(n117[4]), .C1(GND_net), 
          .D1(GND_net), .CIN(n43854), .COUT(n43855), .S0(n21358[2]), 
          .S1(n21358[3]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(108[51:107])
    defparam add_11128_4.INIT0 = 16'h5666;
    defparam add_11128_4.INIT1 = 16'h5666;
    defparam add_11128_4.INJECT1_0 = "NO";
    defparam add_11128_4.INJECT1_1 = "NO";
    CCU2D add_11128_2 (.A0(next_z_linear_velocity_calc_15__N_1577[1]), .B0(next_z_linear_velocity_calc_15__N_1577[2]), 
          .C0(GND_net), .D0(GND_net), .A1(next_z_linear_velocity_calc_15__N_1577[2]), 
          .B1(next_z_linear_velocity_calc_15__N_1577[3]), .C1(GND_net), 
          .D1(GND_net), .COUT(n43854), .S1(n21358[1]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(108[51:107])
    defparam add_11128_2.INIT0 = 16'h7000;
    defparam add_11128_2.INIT1 = 16'h5666;
    defparam add_11128_2.INJECT1_0 = "NO";
    defparam add_11128_2.INJECT1_1 = "NO";
    LUT4 i1_3_lut_adj_280 (.A(\next_state_4__N_1567[2] ), .B(\next_state_4__N_1656[2] ), 
         .C(us_clk_enable_103), .Z(n46653)) /* synthesis lut_function=(A+!((C)+!B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(74[38:48])
    defparam i1_3_lut_adj_280.init = 16'haeae;
    LUT4 i33207_2_lut (.A(next_z_linear_velocity_calc_15__N_1577[1]), .B(n117[3]), 
         .Z(next_z_linear_velocity_calc_15__N_1577[4])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i33207_2_lut.init = 16'h6666;
    LUT4 i20088_2_lut_4_lut (.A(state[2]), .B(state[1]), .C(n52285), .D(sys_clk_enable_252), 
         .Z(n30748)) /* synthesis lut_function=(A (B (D)+!B (C (D)))+!A (D)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(104[17:28])
    defparam i20088_2_lut_4_lut.init = 16'hfd00;
    LUT4 i1_2_lut_rep_497 (.A(state[4]), .B(state[3]), .Z(n52433)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_497.init = 16'heeee;
    LUT4 i1_2_lut_rep_349_3_lut (.A(state[4]), .B(state[3]), .C(state[0]), 
         .Z(n52285)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i1_2_lut_rep_349_3_lut.init = 16'hfefe;
    LUT4 i19_4_lut_3_lut (.A(state[4]), .B(state[3]), .C(state[0]), .Z(n8)) /* synthesis lut_function=(!(A+(B (C)+!B !(C)))) */ ;
    defparam i19_4_lut_3_lut.init = 16'h1414;
    LUT4 i3_4_lut_adj_281 (.A(n52341), .B(n22), .C(n37731), .D(n52342), 
         .Z(n15182)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i3_4_lut_adj_281.init = 16'h0004;
    LUT4 i36_2_lut (.A(\state[2] ), .B(\state[5] ), .Z(n22)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i36_2_lut.init = 16'h6666;
    CCU2D sub_50_add_2_15 (.A0(z_altitude_mm_previous[13]), .B0(z_altitude_mm_latched[13]), 
          .C0(GND_net), .D0(GND_net), .A1(z_altitude_mm_previous[14]), 
          .B1(z_altitude_mm_latched[14]), .C1(GND_net), .D1(GND_net), 
          .CIN(n43841), .S0(n117[13]), .S1(n117[14]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(108[51:99])
    defparam sub_50_add_2_15.INIT0 = 16'h5999;
    defparam sub_50_add_2_15.INIT1 = 16'h5999;
    defparam sub_50_add_2_15.INJECT1_0 = "NO";
    defparam sub_50_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_50_add_2_13 (.A0(z_altitude_mm_previous[11]), .B0(z_altitude_mm_latched[11]), 
          .C0(GND_net), .D0(GND_net), .A1(z_altitude_mm_previous[12]), 
          .B1(z_altitude_mm_latched[12]), .C1(GND_net), .D1(GND_net), 
          .CIN(n43840), .COUT(n43841), .S0(n117[11]), .S1(n117[12]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(108[51:99])
    defparam sub_50_add_2_13.INIT0 = 16'h5999;
    defparam sub_50_add_2_13.INIT1 = 16'h5999;
    defparam sub_50_add_2_13.INJECT1_0 = "NO";
    defparam sub_50_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_50_add_2_11 (.A0(z_altitude_mm_previous[9]), .B0(z_altitude_mm_latched[9]), 
          .C0(GND_net), .D0(GND_net), .A1(z_altitude_mm_previous[10]), 
          .B1(z_altitude_mm_latched[10]), .C1(GND_net), .D1(GND_net), 
          .CIN(n43839), .COUT(n43840), .S0(n117[9]), .S1(n117[10]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(108[51:99])
    defparam sub_50_add_2_11.INIT0 = 16'h5999;
    defparam sub_50_add_2_11.INIT1 = 16'h5999;
    defparam sub_50_add_2_11.INJECT1_0 = "NO";
    defparam sub_50_add_2_11.INJECT1_1 = "NO";
    PFUMX i40920 (.BLUT(n52489), .ALUT(n52490), .C0(state[2]), .Z(next_state_4__N_1576));
    CCU2D sub_50_add_2_9 (.A0(z_altitude_mm_previous[7]), .B0(z_altitude_mm_latched[7]), 
          .C0(GND_net), .D0(GND_net), .A1(z_altitude_mm_previous[8]), 
          .B1(z_altitude_mm_latched[8]), .C1(GND_net), .D1(GND_net), .CIN(n43838), 
          .COUT(n43839), .S0(n117[7]), .S1(n117[8]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(108[51:99])
    defparam sub_50_add_2_9.INIT0 = 16'h5999;
    defparam sub_50_add_2_9.INIT1 = 16'h5999;
    defparam sub_50_add_2_9.INJECT1_0 = "NO";
    defparam sub_50_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_50_add_2_7 (.A0(z_altitude_mm_previous[5]), .B0(z_altitude_mm_latched[5]), 
          .C0(GND_net), .D0(GND_net), .A1(z_altitude_mm_previous[6]), 
          .B1(z_altitude_mm_latched[6]), .C1(GND_net), .D1(GND_net), .CIN(n43837), 
          .COUT(n43838), .S0(n117[5]), .S1(n117[6]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(108[51:99])
    defparam sub_50_add_2_7.INIT0 = 16'h5999;
    defparam sub_50_add_2_7.INIT1 = 16'h5999;
    defparam sub_50_add_2_7.INJECT1_0 = "NO";
    defparam sub_50_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_50_add_2_5 (.A0(z_altitude_mm_previous[3]), .B0(z_altitude_mm_latched[3]), 
          .C0(GND_net), .D0(GND_net), .A1(z_altitude_mm_previous[4]), 
          .B1(z_altitude_mm_latched[4]), .C1(GND_net), .D1(GND_net), .CIN(n43836), 
          .COUT(n43837), .S0(n117[3]), .S1(n117[4]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(108[51:99])
    defparam sub_50_add_2_5.INIT0 = 16'h5999;
    defparam sub_50_add_2_5.INIT1 = 16'h5999;
    defparam sub_50_add_2_5.INJECT1_0 = "NO";
    defparam sub_50_add_2_5.INJECT1_1 = "NO";
    CCU2D sub_50_add_2_3 (.A0(z_altitude_mm_previous[1]), .B0(z_altitude_mm_latched[1]), 
          .C0(GND_net), .D0(GND_net), .A1(z_altitude_mm_previous[2]), 
          .B1(z_altitude_mm_latched[2]), .C1(GND_net), .D1(GND_net), .CIN(n43835), 
          .COUT(n43836), .S0(next_z_linear_velocity_calc_15__N_1577[2]), 
          .S1(next_z_linear_velocity_calc_15__N_1577[3]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(108[51:99])
    defparam sub_50_add_2_3.INIT0 = 16'h5999;
    defparam sub_50_add_2_3.INIT1 = 16'h5999;
    defparam sub_50_add_2_3.INJECT1_0 = "NO";
    defparam sub_50_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_50_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(z_altitude_mm_previous[0]), .B1(z_altitude_mm_latched[0]), 
          .C1(GND_net), .D1(GND_net), .COUT(n43835), .S1(next_z_linear_velocity_calc_15__N_1577[1]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(108[51:99])
    defparam sub_50_add_2_1.INIT0 = 16'h0000;
    defparam sub_50_add_2_1.INIT1 = 16'h5999;
    defparam sub_50_add_2_1.INJECT1_0 = "NO";
    defparam sub_50_add_2_1.INJECT1_1 = "NO";
    LUT4 i32727_4_lut_3_lut_4_lut (.A(\z_linear_velocity[7] ), .B(\z_linear_velocity[4] ), 
         .C(\z_linear_velocity[6] ), .D(\z_linear_velocity[5] ), .Z(n43309)) /* synthesis lut_function=(A (B (D)+!B !((D)+!C))+!A (D)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam i32727_4_lut_3_lut_4_lut.init = 16'hdd20;
    LUT4 i57_2_lut (.A(state[4]), .B(state[0]), .Z(n27)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i57_2_lut.init = 16'h6666;
    FD1P3IX z_linear_velocity_calc_i0_i10 (.D(next_z_linear_velocity_calc_15__N_1577[10]), 
            .SP(sys_clk_enable_257), .CD(n30639), .CK(sys_clk), .Q(\z_linear_velocity[10] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_linear_velocity_calc_i0_i10.GSR = "ENABLED";
    FD1P3IX z_linear_velocity_calc_i0_i11 (.D(next_z_linear_velocity_calc_15__N_1577[11]), 
            .SP(sys_clk_enable_257), .CD(n30639), .CK(sys_clk), .Q(\z_linear_velocity[11] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_linear_velocity_calc_i0_i11.GSR = "ENABLED";
    FD1P3IX z_altitude_mm_latched_i0_i1 (.D(\VL53L1X_range_mm[1] ), .SP(sys_clk_enable_252), 
            .CD(n30748), .CK(sys_clk), .Q(z_altitude_mm_latched[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_altitude_mm_latched_i0_i1.GSR = "ENABLED";
    FD1P3IX z_altitude_mm_latched_i0_i2 (.D(\VL53L1X_range_mm[2] ), .SP(sys_clk_enable_252), 
            .CD(n30748), .CK(sys_clk), .Q(z_altitude_mm_latched[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_altitude_mm_latched_i0_i2.GSR = "ENABLED";
    FD1P3IX z_altitude_mm_latched_i0_i3 (.D(\VL53L1X_range_mm[3] ), .SP(sys_clk_enable_252), 
            .CD(n30748), .CK(sys_clk), .Q(z_altitude_mm_latched[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_altitude_mm_latched_i0_i3.GSR = "ENABLED";
    FD1P3IX z_altitude_mm_latched_i0_i4 (.D(\VL53L1X_range_mm[4] ), .SP(sys_clk_enable_252), 
            .CD(n30748), .CK(sys_clk), .Q(z_altitude_mm_latched[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_altitude_mm_latched_i0_i4.GSR = "ENABLED";
    FD1P3IX z_altitude_mm_latched_i0_i5 (.D(\VL53L1X_range_mm[5] ), .SP(sys_clk_enable_252), 
            .CD(n30748), .CK(sys_clk), .Q(z_altitude_mm_latched[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_altitude_mm_latched_i0_i5.GSR = "ENABLED";
    FD1P3IX z_altitude_mm_latched_i0_i6 (.D(\VL53L1X_range_mm[6] ), .SP(sys_clk_enable_252), 
            .CD(n30748), .CK(sys_clk), .Q(z_altitude_mm_latched[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_altitude_mm_latched_i0_i6.GSR = "ENABLED";
    FD1P3IX z_altitude_mm_latched_i0_i7 (.D(\VL53L1X_range_mm[7] ), .SP(sys_clk_enable_252), 
            .CD(n30748), .CK(sys_clk), .Q(z_altitude_mm_latched[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_altitude_mm_latched_i0_i7.GSR = "ENABLED";
    FD1P3IX z_altitude_mm_latched_i0_i8 (.D(\VL53L1X_range_mm[8] ), .SP(sys_clk_enable_252), 
            .CD(n30748), .CK(sys_clk), .Q(z_altitude_mm_latched[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_altitude_mm_latched_i0_i8.GSR = "ENABLED";
    FD1P3IX z_altitude_mm_latched_i0_i9 (.D(\VL53L1X_range_mm[9] ), .SP(sys_clk_enable_252), 
            .CD(n30748), .CK(sys_clk), .Q(z_altitude_mm_latched[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_altitude_mm_latched_i0_i9.GSR = "ENABLED";
    FD1P3IX z_altitude_mm_latched_i0_i10 (.D(\VL53L1X_range_mm[10] ), .SP(sys_clk_enable_252), 
            .CD(n30748), .CK(sys_clk), .Q(z_altitude_mm_latched[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_altitude_mm_latched_i0_i10.GSR = "ENABLED";
    FD1P3IX z_altitude_mm_latched_i0_i11 (.D(\VL53L1X_range_mm[11] ), .SP(sys_clk_enable_252), 
            .CD(n30748), .CK(sys_clk), .Q(z_altitude_mm_latched[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_altitude_mm_latched_i0_i11.GSR = "ENABLED";
    FD1P3IX z_altitude_mm_latched_i0_i12 (.D(\VL53L1X_range_mm[12] ), .SP(sys_clk_enable_252), 
            .CD(n30748), .CK(sys_clk), .Q(z_altitude_mm_latched[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_altitude_mm_latched_i0_i12.GSR = "ENABLED";
    FD1P3IX z_altitude_mm_latched_i0_i13 (.D(\VL53L1X_range_mm[13] ), .SP(sys_clk_enable_252), 
            .CD(n30748), .CK(sys_clk), .Q(z_altitude_mm_latched[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_altitude_mm_latched_i0_i13.GSR = "ENABLED";
    FD1P3IX z_altitude_mm_latched_i0_i14 (.D(\VL53L1X_range_mm[14] ), .SP(sys_clk_enable_252), 
            .CD(n30748), .CK(sys_clk), .Q(z_altitude_mm_latched[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_altitude_mm_latched_i0_i14.GSR = "ENABLED";
    FD1P3IX z_altitude_mm_previous_i0_i1 (.D(z_altitude_mm_latched[1]), .SP(sys_clk_enable_251), 
            .CD(n30732), .CK(sys_clk), .Q(z_altitude_mm_previous[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_altitude_mm_previous_i0_i1.GSR = "ENABLED";
    FD1P3IX z_altitude_mm_previous_i0_i2 (.D(z_altitude_mm_latched[2]), .SP(sys_clk_enable_251), 
            .CD(n30732), .CK(sys_clk), .Q(z_altitude_mm_previous[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_altitude_mm_previous_i0_i2.GSR = "ENABLED";
    FD1P3IX z_altitude_mm_previous_i0_i3 (.D(z_altitude_mm_latched[3]), .SP(sys_clk_enable_251), 
            .CD(n30732), .CK(sys_clk), .Q(z_altitude_mm_previous[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_altitude_mm_previous_i0_i3.GSR = "ENABLED";
    FD1P3IX z_altitude_mm_previous_i0_i4 (.D(z_altitude_mm_latched[4]), .SP(sys_clk_enable_251), 
            .CD(n30732), .CK(sys_clk), .Q(z_altitude_mm_previous[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_altitude_mm_previous_i0_i4.GSR = "ENABLED";
    FD1P3IX z_altitude_mm_previous_i0_i5 (.D(z_altitude_mm_latched[5]), .SP(sys_clk_enable_251), 
            .CD(n30732), .CK(sys_clk), .Q(z_altitude_mm_previous[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_altitude_mm_previous_i0_i5.GSR = "ENABLED";
    FD1P3IX z_linear_velocity_calc_i0_i12 (.D(next_z_linear_velocity_calc_15__N_1577[12]), 
            .SP(sys_clk_enable_257), .CD(n30639), .CK(sys_clk), .Q(\z_linear_velocity[12] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_linear_velocity_calc_i0_i12.GSR = "ENABLED";
    FD1P3IX z_altitude_mm_previous_i0_i6 (.D(z_altitude_mm_latched[6]), .SP(sys_clk_enable_251), 
            .CD(n30732), .CK(sys_clk), .Q(z_altitude_mm_previous[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_altitude_mm_previous_i0_i6.GSR = "ENABLED";
    FD1P3IX z_altitude_mm_previous_i0_i7 (.D(z_altitude_mm_latched[7]), .SP(sys_clk_enable_251), 
            .CD(n30732), .CK(sys_clk), .Q(z_altitude_mm_previous[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_altitude_mm_previous_i0_i7.GSR = "ENABLED";
    FD1P3IX z_altitude_mm_previous_i0_i8 (.D(z_altitude_mm_latched[8]), .SP(sys_clk_enable_251), 
            .CD(n30732), .CK(sys_clk), .Q(z_altitude_mm_previous[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_altitude_mm_previous_i0_i8.GSR = "ENABLED";
    FD1P3IX z_altitude_mm_previous_i0_i9 (.D(z_altitude_mm_latched[9]), .SP(sys_clk_enable_251), 
            .CD(n30732), .CK(sys_clk), .Q(z_altitude_mm_previous[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_altitude_mm_previous_i0_i9.GSR = "ENABLED";
    FD1P3IX z_altitude_mm_previous_i0_i10 (.D(z_altitude_mm_latched[10]), 
            .SP(sys_clk_enable_251), .CD(n30732), .CK(sys_clk), .Q(z_altitude_mm_previous[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_altitude_mm_previous_i0_i10.GSR = "ENABLED";
    FD1P3IX z_altitude_mm_previous_i0_i11 (.D(z_altitude_mm_latched[11]), 
            .SP(sys_clk_enable_251), .CD(n30732), .CK(sys_clk), .Q(z_altitude_mm_previous[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_altitude_mm_previous_i0_i11.GSR = "ENABLED";
    FD1P3IX z_altitude_mm_previous_i0_i12 (.D(z_altitude_mm_latched[12]), 
            .SP(sys_clk_enable_251), .CD(n30732), .CK(sys_clk), .Q(z_altitude_mm_previous[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_altitude_mm_previous_i0_i12.GSR = "ENABLED";
    FD1P3IX z_altitude_mm_previous_i0_i13 (.D(z_altitude_mm_latched[13]), 
            .SP(sys_clk_enable_251), .CD(n30732), .CK(sys_clk), .Q(z_altitude_mm_previous[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_altitude_mm_previous_i0_i13.GSR = "ENABLED";
    FD1P3IX z_altitude_mm_previous_i0_i14 (.D(z_altitude_mm_latched[14]), 
            .SP(sys_clk_enable_251), .CD(n30732), .CK(sys_clk), .Q(z_altitude_mm_previous[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_altitude_mm_previous_i0_i14.GSR = "ENABLED";
    FD1P3IX z_linear_velocity_calc_i0_i13 (.D(next_z_linear_velocity_calc_15__N_1577[13]), 
            .SP(sys_clk_enable_257), .CD(n30639), .CK(sys_clk), .Q(\z_linear_velocity[13] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_linear_velocity_calc_i0_i13.GSR = "ENABLED";
    FD1P3IX z_linear_velocity_calc_i0_i14 (.D(next_z_linear_velocity_calc_15__N_1577[14]), 
            .SP(sys_clk_enable_257), .CD(n30639), .CK(sys_clk), .Q(\z_linear_velocity[14] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_linear_velocity_calc_i0_i14.GSR = "ENABLED";
    FD1P3IX z_linear_velocity_calc_i0_i15 (.D(next_z_linear_velocity_calc_15__N_1577[15]), 
            .SP(sys_clk_enable_257), .CD(n30639), .CK(sys_clk), .Q(\z_linear_velocity[15] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_linear_velocity_calc_i0_i15.GSR = "ENABLED";
    FD1P3IX z_linear_velocity_calc_i0_i1 (.D(next_z_linear_velocity_calc_15__N_1577[1]), 
            .SP(sys_clk_enable_257), .CD(n30639), .CK(sys_clk), .Q(\z_linear_velocity[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_linear_velocity_calc_i0_i1.GSR = "ENABLED";
    FD1P3IX z_linear_velocity_calc_i0_i2 (.D(next_z_linear_velocity_calc_15__N_1577[2]), 
            .SP(sys_clk_enable_257), .CD(n30639), .CK(sys_clk), .Q(\z_linear_velocity[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_linear_velocity_calc_i0_i2.GSR = "ENABLED";
    FD1P3IX z_linear_velocity_calc_i0_i3 (.D(next_z_linear_velocity_calc_15__N_1577[3]), 
            .SP(sys_clk_enable_257), .CD(n30639), .CK(sys_clk), .Q(\z_linear_velocity[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_linear_velocity_calc_i0_i3.GSR = "ENABLED";
    FD1P3IX z_linear_velocity_calc_i0_i4 (.D(next_z_linear_velocity_calc_15__N_1577[4]), 
            .SP(sys_clk_enable_257), .CD(n30639), .CK(sys_clk), .Q(\z_linear_velocity[4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_linear_velocity_calc_i0_i4.GSR = "ENABLED";
    FD1P3IX z_linear_velocity_calc_i0_i5 (.D(next_z_linear_velocity_calc_15__N_1577[5]), 
            .SP(sys_clk_enable_257), .CD(n30639), .CK(sys_clk), .Q(\z_linear_velocity[5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_linear_velocity_calc_i0_i5.GSR = "ENABLED";
    FD1P3IX z_linear_velocity_calc_i0_i6 (.D(next_z_linear_velocity_calc_15__N_1577[6]), 
            .SP(sys_clk_enable_257), .CD(n30639), .CK(sys_clk), .Q(\z_linear_velocity[6] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_linear_velocity_calc_i0_i6.GSR = "ENABLED";
    FD1P3IX z_linear_velocity_calc_i0_i7 (.D(next_z_linear_velocity_calc_15__N_1577[7]), 
            .SP(sys_clk_enable_257), .CD(n30639), .CK(sys_clk), .Q(\z_linear_velocity[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_linear_velocity_calc_i0_i7.GSR = "ENABLED";
    FD1P3IX z_altitude_mm_previous_i0_i0 (.D(z_altitude_mm_latched[0]), .SP(sys_clk_enable_251), 
            .CD(n30732), .CK(sys_clk), .Q(z_altitude_mm_previous[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_altitude_mm_previous_i0_i0.GSR = "ENABLED";
    FD1P3IX z_altitude_mm_latched_i0_i0 (.D(\VL53L1X_range_mm[0] ), .SP(sys_clk_enable_252), 
            .CD(n30748), .CK(sys_clk), .Q(z_altitude_mm_latched[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_altitude_mm_latched_i0_i0.GSR = "ENABLED";
    FD1P3IX z_linear_velocity_calc_i0_i8 (.D(next_z_linear_velocity_calc_15__N_1577[8]), 
            .SP(sys_clk_enable_257), .CD(n30639), .CK(sys_clk), .Q(\z_linear_velocity[8] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_linear_velocity_calc_i0_i8.GSR = "ENABLED";
    FD1P3IX z_linear_velocity_calc_i0_i9 (.D(next_z_linear_velocity_calc_15__N_1577[9]), 
            .SP(sys_clk_enable_257), .CD(n30639), .CK(sys_clk), .Q(\z_linear_velocity[9] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=28, LSE_RCOL=6, LSE_LLINE=352, LSE_RLINE=358 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/z_linear_velocity_comp.v(58[14] 63[12])
    defparam z_linear_velocity_calc_i0_i9.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module auto_mode_controller
//

module auto_mode_controller (state, resetn_derived_2, count__auto_time_ms_27__N_1647, 
            n53885, us_clk, amc_complete_signal, \amc_debug[0] , next_state_4__N_1666, 
            GND_net, \next_state_14__N_2466[1] , \next_state_4__N_1656[2] , 
            n52214, n4, us_clk_enable_103, \throttle_val[1] , switch_b, 
            \next_auto_state_8__N_1686[7] , \amc_debug[8] , \amc_debug[7] , 
            \amc_debug[6] , \amc_debug[5] , \amc_debug[4] , \amc_debug[3] , 
            \amc_debug[2] , \amc_debug[1] , count__auto_time_ms_27__N_1639, 
            n41683, n41688, n46653, \throttle_val[2] , \throttle_val[3] , 
            \throttle_val[4] , \throttle_val[5] , \throttle_val[6] , \throttle_val[7] , 
            n52213, n48787, n37558, n33315, n52566) /* synthesis syn_module_defined=1 */ ;
    output [4:0]state;
    input resetn_derived_2;
    input count__auto_time_ms_27__N_1647;
    input n53885;
    input us_clk;
    output amc_complete_signal;
    output \amc_debug[0] ;
    input next_state_4__N_1666;
    input GND_net;
    input \next_state_14__N_2466[1] ;
    output \next_state_4__N_1656[2] ;
    input n52214;
    output n4;
    output us_clk_enable_103;
    input \throttle_val[1] ;
    input [1:0]switch_b;
    input \next_auto_state_8__N_1686[7] ;
    output \amc_debug[8] ;
    output \amc_debug[7] ;
    output \amc_debug[6] ;
    output \amc_debug[5] ;
    output \amc_debug[4] ;
    output \amc_debug[3] ;
    output \amc_debug[2] ;
    output \amc_debug[1] ;
    input count__auto_time_ms_27__N_1639;
    output n41683;
    output n41688;
    input n46653;
    input \throttle_val[2] ;
    input \throttle_val[3] ;
    input \throttle_val[4] ;
    input \throttle_val[5] ;
    input \throttle_val[6] ;
    input \throttle_val[7] ;
    output n52213;
    input n48787;
    output n37558;
    output n33315;
    input n52566;
    
    wire next_complete_signal_N_1862 /* synthesis is_clock=1, SET_AS_NETWORK=\AMC/next_complete_signal_N_1862 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(58[9:29])
    wire us_clk /* synthesis SET_AS_NETWORK=us_clk, is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(221[10:16])
    wire next_auto_state_8__N_1765 /* synthesis is_clock=1, SET_AS_NETWORK=\AMC/next_auto_state_8__N_1765 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(76[48:63])
    wire next_state_4__N_1669 /* synthesis is_clock=1, SET_AS_NETWORK=\AMC/next_state_4__N_1669 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(74[38:48])
    
    wire n52313, n48170;
    wire [8:0]auto_state;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(76[36:46])
    wire [8:0]next_auto_state_8__N_1835;
    
    wire n25915, n10, n6, n52310, n52312, n49305, n48672, n88, 
        n52480, n52481, n52482, n30524;
    wire [4:0]next_state;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(74[38:48])
    wire [8:0]next_auto_state;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(76[48:63])
    
    wire next_complete_signal, next_auto_state_8__N_1756, n43822;
    wire [27:0]count__auto_time_ms;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(69[15:34])
    wire [27:0]count__auto_time_ms_27__N_1767;
    
    wire n43823, next_state_4__N_1653, n43821, n52237, n8409, n51604, 
        n8584, n25676, n51603, next_auto_state_8__N_1747, next_auto_state_8__N_1738, 
        next_auto_state_8__N_1729, next_auto_state_8__N_1720, next_auto_state_8__N_1711, 
        next_auto_state_8__N_1702, next_auto_state_8__N_1693, next_auto_state_8__N_1670, 
        n52435, n52571, n52570, n52572, n52426, n52438, n8551, 
        n52198, n52176, n52204, n47375, n30589, n30588, n30586, 
        n30585;
    wire [7:0]throttle_pwm_val_latched;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(64[34:58])
    
    wire n52469, n51, n52308, n8, n4_adj_5179, n48612, n49091, 
        n50694, n50693;
    wire [0:0]n8639;
    
    wire n52191, n12, n4_adj_5180, n7, n8_adj_5181;
    wire [0:0]n8462;
    
    wire n52190, n48049, n30526, n30525, next_auto_state_8__N_1703;
    wire [0:0]n8366;
    
    wire n52189, n43, n48651, n48938, n51605, n4_adj_5182, n91, 
        n52468, n88_adj_5183, n52249, n49361, n52474, n52475, n27592, 
        n44, n30550, n30549, n52325, n34, n30532, n30531, n52326, 
        n52401, n30, n30528;
    wire [27:0]n58;
    
    wire n30534, n30537, n30540, n30543, n30546, n30552, n30555, 
        n30558, n30561, n30564, n30567, us_clk_enable_66, n30570, 
        n30573, n30576, n30579, n30582, n30591, n47358, n48862, 
        n49239, n37959, n30583, n30592, n25, n17, n14, start_flag_N_1875, 
        n48533, n49347, n8_adj_5188, n48795;
    wire [0:0]n8620;
    
    wire n30529, n45_adj_5189, n37_adj_5190, n44_adj_5191, n38_adj_5192, 
        n42_adj_5193, n7_adj_5194, n8_adj_5195, n40_adj_5196, n30541, 
        n30565, n30544, n30574, n30568, n30580, n30538, n30562, 
        n30553, n30535, n30556, n30571, n30577, n30559, n30547, 
        n43834, n43833, n43832, n43831, n19, n24, n14_adj_5197, 
        n22, n16, n43830, n43829, n43828, n43827, n43826, n43825, 
        n43824;
    
    LUT4 i15446_3_lut_4_lut (.A(n52313), .B(n48170), .C(auto_state[7]), 
         .D(next_auto_state_8__N_1835[4]), .Z(n25915)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(159[53:84])
    defparam i15446_3_lut_4_lut.init = 16'hf010;
    PFUMX i22 (.BLUT(n10), .ALUT(n6), .C0(state[4]), .Z(next_complete_signal_N_1862));
    LUT4 i38513_3_lut_4_lut (.A(n52310), .B(n52312), .C(auto_state[2]), 
         .D(auto_state[6]), .Z(n49305)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i38513_3_lut_4_lut.init = 16'hfffe;
    LUT4 i2_3_lut_4_lut (.A(auto_state[5]), .B(n52312), .C(auto_state[3]), 
         .D(auto_state[4]), .Z(n48672)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i2_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_4_lut (.A(auto_state[1]), .B(auto_state[0]), .C(auto_state[2]), 
         .D(auto_state[3]), .Z(n88)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (B (C+(D))+!B (C (D)+!C !(D))))) */ ;
    defparam i1_4_lut_4_lut.init = 16'h0116;
    PFUMX i40914 (.BLUT(n52480), .ALUT(n52481), .C0(auto_state[8]), .Z(n52482));
    LUT4 i1_3_lut_4_lut_4_lut (.A(state[0]), .B(state[1]), .C(state[3]), 
         .D(state[2]), .Z(n10)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (B (C+(D))+!B (C (D)+!C !(D))))) */ ;
    defparam i1_3_lut_4_lut_4_lut.init = 16'h0116;
    FD1S1D i19852 (.D(n53885), .CK(resetn_derived_2), .CD(count__auto_time_ms_27__N_1647), 
           .Q(n30524));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam i19852.GSR = "DISABLED";
    FD1S3AY state_i0 (.D(next_state[0]), .CK(us_clk), .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(123[14] 134[12])
    defparam state_i0.GSR = "ENABLED";
    FD1S3AY auto_state_i0 (.D(next_auto_state[0]), .CK(us_clk), .Q(auto_state[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(123[14] 134[12])
    defparam auto_state_i0.GSR = "ENABLED";
    FD1S3AX complete_signal_386 (.D(next_complete_signal), .CK(us_clk), 
            .Q(amc_complete_signal)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(123[14] 134[12])
    defparam complete_signal_386.GSR = "ENABLED";
    FD1S3AX debug_i1 (.D(auto_state[0]), .CK(us_clk), .Q(\amc_debug[0] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(123[14] 134[12])
    defparam debug_i1.GSR = "ENABLED";
    FD1S1AY next_auto_state_8__I_0_i1 (.D(next_auto_state_8__N_1756), .CK(next_auto_state_8__N_1765), 
            .Q(next_auto_state[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(138[5] 228[8])
    defparam next_auto_state_8__I_0_i1.GSR = "ENABLED";
    FD1S1AY next_state_4__I_50_i1 (.D(next_state_4__N_1666), .CK(next_state_4__N_1669), 
            .Q(next_state[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(138[5] 228[8])
    defparam next_state_4__I_50_i1.GSR = "ENABLED";
    CCU2D sub_8_add_2_5 (.A0(count__auto_time_ms[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count__auto_time_ms[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43822), .COUT(n43823), .S0(count__auto_time_ms_27__N_1767[3]), 
          .S1(count__auto_time_ms_27__N_1767[4]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(90[36:64])
    defparam sub_8_add_2_5.INIT0 = 16'h5555;
    defparam sub_8_add_2_5.INIT1 = 16'h5555;
    defparam sub_8_add_2_5.INJECT1_0 = "NO";
    defparam sub_8_add_2_5.INJECT1_1 = "NO";
    FD1S1A next_complete_signal_I_0 (.D(next_state_4__N_1653), .CK(next_complete_signal_N_1862), 
           .Q(next_complete_signal)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(232[5] 338[8])
    defparam next_complete_signal_I_0.GSR = "ENABLED";
    CCU2D sub_8_add_2_3 (.A0(count__auto_time_ms[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count__auto_time_ms[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43821), .COUT(n43822), .S0(count__auto_time_ms_27__N_1767[1]), 
          .S1(count__auto_time_ms_27__N_1767[2]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(90[36:64])
    defparam sub_8_add_2_3.INIT0 = 16'h5555;
    defparam sub_8_add_2_3.INIT1 = 16'h5555;
    defparam sub_8_add_2_3.INJECT1_0 = "NO";
    defparam sub_8_add_2_3.INJECT1_1 = "NO";
    LUT4 n25915_bdd_4_lut_41338 (.A(n25915), .B(n52237), .C(n8409), .D(auto_state[5]), 
         .Z(n51604)) /* synthesis lut_function=(A ((C+!(D))+!B)+!A (B (C)+!B (C+(D)))) */ ;
    defparam n25915_bdd_4_lut_41338.init = 16'hf3fa;
    LUT4 n25915_bdd_4_lut_40542 (.A(n52237), .B(n8584), .C(n25676), .D(auto_state[0]), 
         .Z(n51603)) /* synthesis lut_function=((B (C)+!B (D))+!A) */ ;
    defparam n25915_bdd_4_lut_40542.init = 16'hf7d5;
    FD1S1A next_auto_state_8__I_0_i2 (.D(next_auto_state_8__N_1747), .CK(next_auto_state_8__N_1765), 
           .Q(next_auto_state[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(138[5] 228[8])
    defparam next_auto_state_8__I_0_i2.GSR = "ENABLED";
    FD1S1A next_auto_state_8__I_0_i3 (.D(next_auto_state_8__N_1738), .CK(next_auto_state_8__N_1765), 
           .Q(next_auto_state[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(138[5] 228[8])
    defparam next_auto_state_8__I_0_i3.GSR = "ENABLED";
    FD1S1A next_auto_state_8__I_0_i4 (.D(next_auto_state_8__N_1729), .CK(next_auto_state_8__N_1765), 
           .Q(next_auto_state[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(138[5] 228[8])
    defparam next_auto_state_8__I_0_i4.GSR = "ENABLED";
    FD1S1A next_auto_state_8__I_0_i5 (.D(next_auto_state_8__N_1720), .CK(next_auto_state_8__N_1765), 
           .Q(next_auto_state[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(138[5] 228[8])
    defparam next_auto_state_8__I_0_i5.GSR = "ENABLED";
    FD1S1A next_auto_state_8__I_0_i6 (.D(next_auto_state_8__N_1711), .CK(next_auto_state_8__N_1765), 
           .Q(next_auto_state[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(138[5] 228[8])
    defparam next_auto_state_8__I_0_i6.GSR = "ENABLED";
    FD1S1A next_auto_state_8__I_0_i7 (.D(next_auto_state_8__N_1702), .CK(next_auto_state_8__N_1765), 
           .Q(next_auto_state[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(138[5] 228[8])
    defparam next_auto_state_8__I_0_i7.GSR = "ENABLED";
    FD1S1A next_auto_state_8__I_0_i8 (.D(next_auto_state_8__N_1693), .CK(next_auto_state_8__N_1765), 
           .Q(next_auto_state[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(138[5] 228[8])
    defparam next_auto_state_8__I_0_i8.GSR = "ENABLED";
    FD1S1A next_auto_state_8__I_0_i9 (.D(next_auto_state_8__N_1670), .CK(next_auto_state_8__N_1765), 
           .Q(next_auto_state[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(138[5] 228[8])
    defparam next_auto_state_8__I_0_i9.GSR = "ENABLED";
    LUT4 mux_3820_i2_3_lut_4_lut_4_lut_then_4_lut (.A(n52435), .B(\next_state_14__N_2466[1] ), 
         .C(state[4]), .D(state[1]), .Z(n52571)) /* synthesis lut_function=(!(A+!(B+(C+(D))))) */ ;
    defparam mux_3820_i2_3_lut_4_lut_4_lut_then_4_lut.init = 16'h5554;
    LUT4 mux_3820_i2_3_lut_4_lut_4_lut_else_4_lut (.A(n52435), .B(\next_state_4__N_1656[2] ), 
         .C(state[4]), .D(state[1]), .Z(n52570)) /* synthesis lut_function=(!(A+!((C+!(D))+!B))) */ ;
    defparam mux_3820_i2_3_lut_4_lut_4_lut_else_4_lut.init = 16'h5155;
    FD1S1I next_state_4__I_50_i2 (.D(n52572), .CK(next_state_4__N_1669), 
           .CD(n52214), .Q(next_state[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(138[5] 228[8])
    defparam next_state_4__I_50_i2.GSR = "ENABLED";
    CCU2D sub_8_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(n52426), .B1(GND_net), .C1(GND_net), .D1(GND_net), .COUT(n43821), 
          .S1(count__auto_time_ms_27__N_1767[0]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(90[36:64])
    defparam sub_8_add_2_1.INIT0 = 16'hF000;
    defparam sub_8_add_2_1.INIT1 = 16'h5555;
    defparam sub_8_add_2_1.INJECT1_0 = "NO";
    defparam sub_8_add_2_1.INJECT1_1 = "NO";
    LUT4 i47_2_lut_rep_502 (.A(state[0]), .B(state[1]), .Z(n52438)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(254[13] 282[20])
    defparam i47_2_lut_rep_502.init = 16'h6666;
    LUT4 i6402_2_lut_rep_240_3_lut (.A(n8551), .B(n52198), .C(n8409), 
         .Z(n52176)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(157[17] 224[24])
    defparam i6402_2_lut_rep_240_3_lut.init = 16'hfbfb;
    LUT4 i3_3_lut_4_lut (.A(n8551), .B(n52198), .C(n52204), .D(n8584), 
         .Z(n47375)) /* synthesis lut_function=(A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(157[17] 224[24])
    defparam i3_3_lut_4_lut.init = 16'h8000;
    LUT4 i19918_3_lut (.A(n30589), .B(n30588), .C(n30524), .Z(count__auto_time_ms[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam i19918_3_lut.init = 16'hcaca;
    LUT4 i19915_3_lut (.A(n30586), .B(n30585), .C(n30524), .Z(count__auto_time_ms[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam i19915_3_lut.init = 16'hcaca;
    LUT4 state_2__bdd_4_lut (.A(state[2]), .B(state[3]), .C(state[4]), 
         .D(state[1]), .Z(n4)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+(C (D)+!C !(D)))) */ ;
    defparam state_2__bdd_4_lut.init = 16'hfeed;
    FD1P3AX throttle_pwm_val_latched__i1 (.D(\throttle_val[1] ), .SP(us_clk_enable_103), 
            .CK(us_clk), .Q(throttle_pwm_val_latched[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(123[14] 134[12])
    defparam throttle_pwm_val_latched__i1.GSR = "ENABLED";
    LUT4 i1_4_lut_then_4_lut (.A(state[1]), .B(state[2]), .C(state[3]), 
         .D(state[4]), .Z(n52469)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(254[13] 282[20])
    defparam i1_4_lut_then_4_lut.init = 16'h0001;
    LUT4 i39846_2_lut_3_lut_4_lut (.A(n52438), .B(n52435), .C(n52214), 
         .D(state[4]), .Z(n51)) /* synthesis lut_function=(!(A (B (C)+!B (C+!(D)))+!A (C))) */ ;
    defparam i39846_2_lut_3_lut_4_lut.init = 16'h0f0d;
    LUT4 i2_4_lut (.A(n52308), .B(n8), .C(n4_adj_5179), .D(n48612), 
         .Z(next_auto_state_8__N_1765)) /* synthesis lut_function=(A ((D)+!B)+!A ((C+(D))+!B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(156[18] 225[16])
    defparam i2_4_lut.init = 16'hff73;
    LUT4 i1_4_lut (.A(n49091), .B(auto_state[4]), .C(n50694), .D(auto_state[5]), 
         .Z(n4_adj_5179)) /* synthesis lut_function=(!(A (B+(D))+!A (B+((D)+!C)))) */ ;
    defparam i1_4_lut.init = 16'h0032;
    LUT4 auto_state_6__bdd_4_lut_39988 (.A(auto_state[7]), .B(auto_state[8]), 
         .C(auto_state[1]), .D(auto_state[0]), .Z(n50693)) /* synthesis lut_function=(!(A+(B (C+(D))+!B (C (D)+!C !(D))))) */ ;
    defparam auto_state_6__bdd_4_lut_39988.init = 16'h0114;
    LUT4 n50693_bdd_2_lut (.A(n50693), .B(auto_state[6]), .Z(n50694)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam n50693_bdd_2_lut.init = 16'h2222;
    LUT4 next_auto_state_8__I_61_4_lut (.A(n8639[0]), .B(auto_state[1]), 
         .C(n8), .D(n52191), .Z(next_auto_state_8__N_1747)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(156[18] 225[16])
    defparam next_auto_state_8__I_61_4_lut.init = 16'hac0c;
    LUT4 i21080_4_lut (.A(auto_state[1]), .B(auto_state[2]), .C(n8), .D(n47375), 
         .Z(next_auto_state_8__N_1738)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B ((D)+!C)+!B (C (D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(76[48:63])
    defparam i21080_4_lut.init = 16'h5c0c;
    LUT4 i3_4_lut (.A(auto_state[6]), .B(n48672), .C(n12), .D(auto_state[0]), 
         .Z(n8584)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i3_4_lut.init = 16'h0010;
    LUT4 i19_2_lut (.A(auto_state[2]), .B(auto_state[1]), .Z(n12)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(76[36:46])
    defparam i19_2_lut.init = 16'h6666;
    LUT4 i21076_4_lut (.A(n47375), .B(auto_state[3]), .C(n8), .D(n4_adj_5180), 
         .Z(next_auto_state_8__N_1729)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(76[48:63])
    defparam i21076_4_lut.init = 16'hac0c;
    LUT4 i1_2_lut (.A(switch_b[0]), .B(auto_state[1]), .Z(n4_adj_5180)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(123[14] 134[12])
    defparam i1_2_lut.init = 16'h8888;
    LUT4 i21111_4_lut (.A(n7), .B(auto_state[4]), .C(n8), .D(n8_adj_5181), 
         .Z(next_auto_state_8__N_1720)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(76[48:63])
    defparam i21111_4_lut.init = 16'hac0c;
    LUT4 i101_2_lut (.A(\next_auto_state_8__N_1686[7] ), .B(switch_b[1]), 
         .Z(next_auto_state_8__N_1835[4])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(211[58:110])
    defparam i101_2_lut.init = 16'h8888;
    LUT4 next_auto_state_8__I_57_4_lut (.A(n8462[0]), .B(auto_state[5]), 
         .C(n8), .D(n52190), .Z(next_auto_state_8__N_1711)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((C)+!B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(156[18] 225[16])
    defparam next_auto_state_8__I_57_4_lut.init = 16'h0cac;
    LUT4 mux_3963_i1_4_lut (.A(auto_state[5]), .B(auto_state[3]), .C(n8409), 
         .D(n48049), .Z(n8462[0])) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(157[17] 224[24])
    defparam mux_3963_i1_4_lut.init = 16'hcac0;
    LUT4 i19855_3_lut (.A(n30526), .B(n30525), .C(n30524), .Z(count__auto_time_ms[27])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam i19855_3_lut.init = 16'hcaca;
    LUT4 next_auto_state_8__I_56_3_lut (.A(next_auto_state_8__N_1703), .B(auto_state[6]), 
         .C(n8), .Z(next_auto_state_8__N_1702)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(156[18] 225[16])
    defparam next_auto_state_8__I_56_3_lut.init = 16'hacac;
    LUT4 next_auto_state_8__I_55_4_lut (.A(n8366[0]), .B(auto_state[7]), 
         .C(n8), .D(n52176), .Z(next_auto_state_8__N_1693)) /* synthesis lut_function=(!(A (B (C (D))+!B ((D)+!C))+!A ((C)+!B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(156[18] 225[16])
    defparam next_auto_state_8__I_55_4_lut.init = 16'h0cac;
    LUT4 mux_3889_i1_4_lut (.A(\next_auto_state_8__N_1686[7] ), .B(n52189), 
         .C(auto_state[5]), .D(n25915), .Z(n8366[0])) /* synthesis lut_function=(A (B (C+!(D))+!B !(C+(D)))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(157[17] 224[24])
    defparam mux_3889_i1_4_lut.init = 16'hc0ca;
    LUT4 i3_4_lut_adj_255 (.A(auto_state[0]), .B(n48049), .C(n8584), .D(n43), 
         .Z(n48651)) /* synthesis lut_function=(!(A+((C+!(D))+!B))) */ ;
    defparam i3_4_lut_adj_255.init = 16'h0400;
    LUT4 i2_3_lut (.A(n52198), .B(n8409), .C(auto_state[3]), .Z(n48938)) /* synthesis lut_function=(!(((C)+!B)+!A)) */ ;
    defparam i2_3_lut.init = 16'h0808;
    LUT4 i1_2_lut_rep_372 (.A(auto_state[3]), .B(auto_state[2]), .Z(n52308)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_372.init = 16'heeee;
    LUT4 next_auto_state_8__I_52_4_lut (.A(n51605), .B(auto_state[8]), .C(n8), 
         .D(n4_adj_5182), .Z(next_auto_state_8__N_1670)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B (C (D))+!B ((D)+!C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(156[18] 225[16])
    defparam next_auto_state_8__I_52_4_lut.init = 16'h0c5c;
    LUT4 i2_3_lut_4_lut_adj_256 (.A(auto_state[3]), .B(auto_state[2]), .C(auto_state[5]), 
         .D(auto_state[4]), .Z(n91)) /* synthesis lut_function=(!(A+(B+(C (D)+!C !(D))))) */ ;
    defparam i2_3_lut_4_lut_adj_256.init = 16'h0110;
    LUT4 i1_4_lut_else_4_lut (.A(state[1]), .B(state[2]), .C(state[3]), 
         .D(state[4]), .Z(n52468)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (B (C+(D))+!B (C (D)+!C !(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(254[13] 282[20])
    defparam i1_4_lut_else_4_lut.init = 16'h0116;
    LUT4 i2_3_lut_4_lut_adj_257 (.A(auto_state[2]), .B(auto_state[3]), .C(auto_state[5]), 
         .D(auto_state[4]), .Z(n88_adj_5183)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A ((C+(D))+!B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(76[36:46])
    defparam i2_3_lut_4_lut_adj_257.init = 16'h0006;
    LUT4 i25745_2_lut_rep_374 (.A(auto_state[0]), .B(auto_state[1]), .Z(n52310)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i25745_2_lut_rep_374.init = 16'heeee;
    LUT4 i25876_2_lut_rep_376 (.A(auto_state[8]), .B(auto_state[7]), .Z(n52312)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i25876_2_lut_rep_376.init = 16'heeee;
    LUT4 i2_4_lut_adj_258 (.A(n88_adj_5183), .B(n52249), .C(n91), .D(auto_state[6]), 
         .Z(n48612)) /* synthesis lut_function=(!(A (B+(D))+!A (B+((D)+!C)))) */ ;
    defparam i2_4_lut_adj_258.init = 16'h0032;
    LUT4 i38566_2_lut_3_lut (.A(auto_state[8]), .B(auto_state[7]), .C(auto_state[6]), 
         .Z(n49361)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i38566_2_lut_3_lut.init = 16'hfefe;
    LUT4 i37570_2_lut_rep_313_3_lut_4_lut (.A(auto_state[8]), .B(auto_state[7]), 
         .C(auto_state[1]), .D(auto_state[0]), .Z(n52249)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i37570_2_lut_rep_313_3_lut_4_lut.init = 16'hfffe;
    LUT4 i12143_2_lut_rep_377 (.A(throttle_pwm_val_latched[6]), .B(throttle_pwm_val_latched[7]), 
         .Z(n52313)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(159[53:84])
    defparam i12143_2_lut_rep_377.init = 16'heeee;
    LUT4 i2_2_lut_3_lut_4_lut (.A(throttle_pwm_val_latched[6]), .B(throttle_pwm_val_latched[7]), 
         .C(auto_state[7]), .D(n48170), .Z(n7)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(159[53:84])
    defparam i2_2_lut_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i2_2_lut_rep_268_3_lut_4_lut (.A(throttle_pwm_val_latched[6]), .B(throttle_pwm_val_latched[7]), 
         .C(\next_auto_state_8__N_1686[7] ), .D(n48170), .Z(n52204)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(159[53:84])
    defparam i2_2_lut_rep_268_3_lut_4_lut.init = 16'hf0e0;
    LUT4 i1_2_lut_rep_301_3_lut (.A(throttle_pwm_val_latched[6]), .B(throttle_pwm_val_latched[7]), 
         .C(n48170), .Z(n52237)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(159[53:84])
    defparam i1_2_lut_rep_301_3_lut.init = 16'hfefe;
    LUT4 i1_4_lut_then_4_lut_adj_259 (.A(auto_state[5]), .B(auto_state[6]), 
         .C(auto_state[4]), .D(auto_state[7]), .Z(n52481)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i1_4_lut_then_4_lut_adj_259.init = 16'h0001;
    PFUMX i40910 (.BLUT(n52474), .ALUT(n52475), .C0(auto_state[6]), .Z(n8551));
    LUT4 i1_3_lut_rep_262 (.A(auto_state[0]), .B(n27592), .C(n44), .Z(n52198)) /* synthesis lut_function=(A (B)+!A (B+(C))) */ ;
    defparam i1_3_lut_rep_262.init = 16'hdcdc;
    LUT4 i2_4_lut_adj_260 (.A(auto_state[8]), .B(auto_state[6]), .C(n52310), 
         .D(auto_state[7]), .Z(n49091)) /* synthesis lut_function=(!(A+(B (C+(D))+!B (C+!(D))))) */ ;
    defparam i2_4_lut_adj_260.init = 16'h0104;
    LUT4 i6370_2_lut_rep_255_4_lut (.A(auto_state[0]), .B(n27592), .C(n44), 
         .D(n8551), .Z(n52191)) /* synthesis lut_function=(A (B (D))+!A (B (D)+!B (C (D)))) */ ;
    defparam i6370_2_lut_rep_255_4_lut.init = 16'hdc00;
    LUT4 i1_2_lut_adj_261 (.A(n44), .B(n27592), .Z(n43)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_adj_261.init = 16'heeee;
    LUT4 i19879_3_lut_rep_389 (.A(n30550), .B(n30549), .C(n30524), .Z(n52325)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam i19879_3_lut_rep_389.init = 16'hcaca;
    LUT4 i10_2_lut_4_lut (.A(n30550), .B(n30549), .C(n30524), .D(count__auto_time_ms[7]), 
         .Z(n34)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam i10_2_lut_4_lut.init = 16'hca00;
    LUT4 i6399_2_lut_rep_254_4_lut (.A(auto_state[0]), .B(n27592), .C(n44), 
         .D(n8551), .Z(n52190)) /* synthesis lut_function=(A ((D)+!B)+!A (B (D)+!B ((D)+!C))) */ ;
    defparam i6399_2_lut_rep_254_4_lut.init = 16'hff23;
    LUT4 i19861_3_lut_rep_390 (.A(n30532), .B(n30531), .C(n30524), .Z(n52326)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam i19861_3_lut_rep_390.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut (.A(auto_state[0]), .B(n27592), .C(n44), .D(\next_auto_state_8__N_1686[7] ), 
         .Z(n4_adj_5182)) /* synthesis lut_function=(A ((D)+!B)+!A (B (D)+!B ((D)+!C))) */ ;
    defparam i1_2_lut_4_lut.init = 16'hff23;
    LUT4 i1_2_lut_rep_465 (.A(auto_state[1]), .B(\next_auto_state_8__N_1686[7] ), 
         .Z(n52401)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(123[14] 134[12])
    defparam i1_2_lut_rep_465.init = 16'h8888;
    LUT4 i6_2_lut_4_lut (.A(n30532), .B(n30531), .C(n30524), .D(count__auto_time_ms[2]), 
         .Z(n30)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam i6_2_lut_4_lut.init = 16'hca00;
    LUT4 i1_2_lut_3_lut (.A(auto_state[1]), .B(\next_auto_state_8__N_1686[7] ), 
         .C(switch_b[0]), .Z(n25676)) /* synthesis lut_function=(A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(123[14] 134[12])
    defparam i1_2_lut_3_lut.init = 16'h8080;
    FD1S3AX debug_i9 (.D(auto_state[8]), .CK(us_clk), .Q(\amc_debug[8] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(123[14] 134[12])
    defparam debug_i9.GSR = "ENABLED";
    FD1S3AX debug_i8 (.D(auto_state[7]), .CK(us_clk), .Q(\amc_debug[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(123[14] 134[12])
    defparam debug_i8.GSR = "ENABLED";
    FD1S3AX debug_i7 (.D(auto_state[6]), .CK(us_clk), .Q(\amc_debug[6] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(123[14] 134[12])
    defparam debug_i7.GSR = "ENABLED";
    FD1S3AX debug_i6 (.D(auto_state[5]), .CK(us_clk), .Q(\amc_debug[5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(123[14] 134[12])
    defparam debug_i6.GSR = "ENABLED";
    FD1S3AX debug_i5 (.D(auto_state[4]), .CK(us_clk), .Q(\amc_debug[4] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(123[14] 134[12])
    defparam debug_i5.GSR = "ENABLED";
    FD1S3AX debug_i4 (.D(auto_state[3]), .CK(us_clk), .Q(\amc_debug[3] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(123[14] 134[12])
    defparam debug_i4.GSR = "ENABLED";
    FD1S3AX debug_i3 (.D(auto_state[2]), .CK(us_clk), .Q(\amc_debug[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(123[14] 134[12])
    defparam debug_i3.GSR = "ENABLED";
    FD1S3AX debug_i2 (.D(auto_state[1]), .CK(us_clk), .Q(\amc_debug[1] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(123[14] 134[12])
    defparam debug_i2.GSR = "ENABLED";
    FD1S3AX auto_state_i8 (.D(next_auto_state[8]), .CK(us_clk), .Q(auto_state[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(123[14] 134[12])
    defparam auto_state_i8.GSR = "ENABLED";
    FD1S3AX auto_state_i7 (.D(next_auto_state[7]), .CK(us_clk), .Q(auto_state[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(123[14] 134[12])
    defparam auto_state_i7.GSR = "ENABLED";
    FD1S3AX auto_state_i6 (.D(next_auto_state[6]), .CK(us_clk), .Q(auto_state[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(123[14] 134[12])
    defparam auto_state_i6.GSR = "ENABLED";
    FD1S3AX auto_state_i5 (.D(next_auto_state[5]), .CK(us_clk), .Q(auto_state[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(123[14] 134[12])
    defparam auto_state_i5.GSR = "ENABLED";
    FD1S3AX auto_state_i4 (.D(next_auto_state[4]), .CK(us_clk), .Q(auto_state[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(123[14] 134[12])
    defparam auto_state_i4.GSR = "ENABLED";
    FD1S3AX auto_state_i3 (.D(next_auto_state[3]), .CK(us_clk), .Q(auto_state[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(123[14] 134[12])
    defparam auto_state_i3.GSR = "ENABLED";
    FD1S3AX auto_state_i2 (.D(next_auto_state[2]), .CK(us_clk), .Q(auto_state[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(123[14] 134[12])
    defparam auto_state_i2.GSR = "ENABLED";
    FD1S3AX auto_state_i1 (.D(next_auto_state[1]), .CK(us_clk), .Q(auto_state[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(123[14] 134[12])
    defparam auto_state_i1.GSR = "ENABLED";
    FD1S3AX state_i4 (.D(next_state[4]), .CK(us_clk), .Q(state[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(123[14] 134[12])
    defparam state_i4.GSR = "ENABLED";
    FD1S3AX state_i3 (.D(next_state[3]), .CK(us_clk), .Q(state[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(123[14] 134[12])
    defparam state_i3.GSR = "ENABLED";
    FD1S3AX state_i2 (.D(next_state[2]), .CK(us_clk), .Q(state[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(123[14] 134[12])
    defparam state_i2.GSR = "ENABLED";
    FD1S3AX state_i1 (.D(next_state[1]), .CK(us_clk), .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(123[14] 134[12])
    defparam state_i1.GSR = "ENABLED";
    FD1S3AY count__auto_time_ms_i0_i26_19856_19857_set (.D(n58[26]), .CK(us_clk), 
            .Q(n30528)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i26_19856_19857_set.GSR = "ENABLED";
    FD1S3AY count__auto_time_ms_i0_i25_19859_19860_set (.D(n58[25]), .CK(us_clk), 
            .Q(n30531)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i25_19859_19860_set.GSR = "ENABLED";
    FD1S3AY count__auto_time_ms_i0_i24_19862_19863_set (.D(n58[24]), .CK(us_clk), 
            .Q(n30534)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i24_19862_19863_set.GSR = "ENABLED";
    FD1S3AY count__auto_time_ms_i0_i23_19865_19866_set (.D(n58[23]), .CK(us_clk), 
            .Q(n30537)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i23_19865_19866_set.GSR = "ENABLED";
    FD1S3AY count__auto_time_ms_i0_i22_19868_19869_set (.D(n58[22]), .CK(us_clk), 
            .Q(n30540)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i22_19868_19869_set.GSR = "ENABLED";
    FD1S3AY count__auto_time_ms_i0_i21_19871_19872_set (.D(n58[21]), .CK(us_clk), 
            .Q(n30543)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i21_19871_19872_set.GSR = "ENABLED";
    FD1S3AY count__auto_time_ms_i0_i20_19874_19875_set (.D(n58[20]), .CK(us_clk), 
            .Q(n30546)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i20_19874_19875_set.GSR = "ENABLED";
    FD1S3AY count__auto_time_ms_i0_i19_19877_19878_set (.D(n58[19]), .CK(us_clk), 
            .Q(n30549)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i19_19877_19878_set.GSR = "ENABLED";
    FD1S3AY count__auto_time_ms_i0_i18_19880_19881_set (.D(n58[18]), .CK(us_clk), 
            .Q(n30552)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i18_19880_19881_set.GSR = "ENABLED";
    FD1S3AY count__auto_time_ms_i0_i17_19883_19884_set (.D(n58[17]), .CK(us_clk), 
            .Q(n30555)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i17_19883_19884_set.GSR = "ENABLED";
    FD1S3AY count__auto_time_ms_i0_i16_19886_19887_set (.D(n58[16]), .CK(us_clk), 
            .Q(n30558)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i16_19886_19887_set.GSR = "ENABLED";
    FD1S3AY count__auto_time_ms_i0_i15_19889_19890_set (.D(n58[15]), .CK(us_clk), 
            .Q(n30561)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i15_19889_19890_set.GSR = "ENABLED";
    FD1S3AY count__auto_time_ms_i0_i14_19892_19893_set (.D(n58[14]), .CK(us_clk), 
            .Q(n30564)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i14_19892_19893_set.GSR = "ENABLED";
    FD1S3AY count__auto_time_ms_i0_i12_19895_19896_set (.D(n58[12]), .CK(us_clk), 
            .Q(n30567)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i12_19895_19896_set.GSR = "ENABLED";
    FD1P3BX count__auto_time_ms_i0_i13 (.D(count__auto_time_ms_27__N_1767[13]), 
            .SP(us_clk_enable_66), .CK(us_clk), .PD(count__auto_time_ms_27__N_1639), 
            .Q(count__auto_time_ms[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i13.GSR = "DISABLED";
    FD1S3AY count__auto_time_ms_i0_i11_19898_19899_set (.D(n58[11]), .CK(us_clk), 
            .Q(n30570)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i11_19898_19899_set.GSR = "ENABLED";
    FD1S3AY count__auto_time_ms_i0_i7_19901_19902_set (.D(n58[7]), .CK(us_clk), 
            .Q(n30573)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i7_19901_19902_set.GSR = "ENABLED";
    FD1P3BX count__auto_time_ms_i0_i10 (.D(count__auto_time_ms_27__N_1767[10]), 
            .SP(us_clk_enable_66), .CK(us_clk), .PD(count__auto_time_ms_27__N_1639), 
            .Q(count__auto_time_ms[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i10.GSR = "DISABLED";
    FD1P3BX count__auto_time_ms_i0_i9 (.D(count__auto_time_ms_27__N_1767[9]), 
            .SP(us_clk_enable_66), .CK(us_clk), .PD(count__auto_time_ms_27__N_1639), 
            .Q(count__auto_time_ms[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i9.GSR = "DISABLED";
    FD1P3BX count__auto_time_ms_i0_i8 (.D(count__auto_time_ms_27__N_1767[8]), 
            .SP(us_clk_enable_66), .CK(us_clk), .PD(count__auto_time_ms_27__N_1639), 
            .Q(count__auto_time_ms[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i8.GSR = "DISABLED";
    FD1S3AY count__auto_time_ms_i0_i6_19904_19905_set (.D(n58[6]), .CK(us_clk), 
            .Q(n30576)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i6_19904_19905_set.GSR = "ENABLED";
    FD1S3AY count__auto_time_ms_i0_i5_19907_19908_set (.D(n58[5]), .CK(us_clk), 
            .Q(n30579)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i5_19907_19908_set.GSR = "ENABLED";
    FD1S3AY count__auto_time_ms_i0_i3_19910_19911_set (.D(n58[3]), .CK(us_clk), 
            .Q(n30582)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i3_19910_19911_set.GSR = "ENABLED";
    FD1P3BX count__auto_time_ms_i0_i4 (.D(count__auto_time_ms_27__N_1767[4]), 
            .SP(us_clk_enable_66), .CK(us_clk), .PD(count__auto_time_ms_27__N_1639), 
            .Q(count__auto_time_ms[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i4.GSR = "DISABLED";
    FD1S3AY count__auto_time_ms_i0_i2_19913_19914_set (.D(n58[2]), .CK(us_clk), 
            .Q(n30585)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i2_19913_19914_set.GSR = "ENABLED";
    FD1S3AY count__auto_time_ms_i0_i1_19916_19917_set (.D(n58[1]), .CK(us_clk), 
            .Q(n30588)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i1_19916_19917_set.GSR = "ENABLED";
    FD1S3AY count__auto_time_ms_i0_i0_19919_19920_set (.D(n58[0]), .CK(us_clk), 
            .Q(n30591)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i0_19919_19920_set.GSR = "ENABLED";
    LUT4 i1_2_lut_3_lut_4_lut (.A(n52313), .B(n48170), .C(count__auto_time_ms[27]), 
         .D(\next_auto_state_8__N_1686[7] ), .Z(n48049)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(159[53:84])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0e00;
    LUT4 i39666_3_lut (.A(state[4]), .B(n47358), .C(state[2]), .Z(us_clk_enable_103)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(277[17:31])
    defparam i39666_3_lut.init = 16'h1010;
    LUT4 i1_2_lut_adj_262 (.A(\amc_debug[7] ), .B(\amc_debug[4] ), .Z(n41683)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(123[14] 134[12])
    defparam i1_2_lut_adj_262.init = 16'hdddd;
    LUT4 i1_2_lut_adj_263 (.A(\amc_debug[0] ), .B(\amc_debug[3] ), .Z(n41688)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(123[14] 134[12])
    defparam i1_2_lut_adj_263.init = 16'hbbbb;
    LUT4 next_auto_state_8__I_62_3_lut (.A(n48862), .B(auto_state[0]), .C(n8), 
         .Z(next_auto_state_8__N_1756)) /* synthesis lut_function=(!(A ((C)+!B)+!A !(B+(C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(156[18] 225[16])
    defparam next_auto_state_8__I_62_3_lut.init = 16'h5c5c;
    LUT4 i2_4_lut_adj_264 (.A(n49239), .B(n48170), .C(n52313), .D(n52198), 
         .Z(n48862)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;
    defparam i2_4_lut_adj_264.init = 16'hfeff;
    FD1S3AX start_flag_383 (.D(n46653), .CK(us_clk), .Q(\next_state_4__N_1656[2] )) /* synthesis lse_init_val=0, LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(98[14] 105[42])
    defparam start_flag_383.GSR = "ENABLED";
    LUT4 i38449_4_lut (.A(n8551), .B(n8409), .C(auto_state[7]), .D(auto_state[5]), 
         .Z(n49239)) /* synthesis lut_function=(!(A+!(B+!(C+(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(157[17] 224[24])
    defparam i38449_4_lut.init = 16'h4445;
    LUT4 i2_4_lut_adj_265 (.A(throttle_pwm_val_latched[4]), .B(n37959), 
         .C(throttle_pwm_val_latched[5]), .D(throttle_pwm_val_latched[3]), 
         .Z(n48170)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(159[53:84])
    defparam i2_4_lut_adj_265.init = 16'hfefa;
    LUT4 i1_4_lut_then_4_lut_adj_266 (.A(n48672), .B(auto_state[0]), .C(auto_state[1]), 
         .D(auto_state[2]), .Z(n52475)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i1_4_lut_then_4_lut_adj_266.init = 16'h0001;
    LUT4 i27282_2_lut (.A(throttle_pwm_val_latched[1]), .B(throttle_pwm_val_latched[2]), 
         .Z(n37959)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i27282_2_lut.init = 16'heeee;
    LUT4 i3_4_lut_adj_267 (.A(n88), .B(n49361), .C(auto_state[4]), .D(auto_state[5]), 
         .Z(n27592)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i3_4_lut_adj_267.init = 16'h0002;
    LUT4 i1_4_lut_else_4_lut_adj_268 (.A(n48672), .B(auto_state[0]), .C(auto_state[1]), 
         .D(auto_state[2]), .Z(n52474)) /* synthesis lut_function=(!(A+(B (C+(D))+!B (C (D)+!C !(D))))) */ ;
    defparam i1_4_lut_else_4_lut_adj_268.init = 16'h0114;
    LUT4 i3_3_lut_4_lut_adj_269 (.A(n8409), .B(n52190), .C(auto_state[5]), 
         .D(next_auto_state_8__N_1835[4]), .Z(n8_adj_5181)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(157[17] 224[24])
    defparam i3_3_lut_4_lut_adj_269.init = 16'h0100;
    FD1P3AX throttle_pwm_val_latched__i2 (.D(\throttle_val[2] ), .SP(us_clk_enable_103), 
            .CK(us_clk), .Q(throttle_pwm_val_latched[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(123[14] 134[12])
    defparam throttle_pwm_val_latched__i2.GSR = "ENABLED";
    FD1P3AX throttle_pwm_val_latched__i3 (.D(\throttle_val[3] ), .SP(us_clk_enable_103), 
            .CK(us_clk), .Q(throttle_pwm_val_latched[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(123[14] 134[12])
    defparam throttle_pwm_val_latched__i3.GSR = "ENABLED";
    FD1P3AX throttle_pwm_val_latched__i4 (.D(\throttle_val[4] ), .SP(us_clk_enable_103), 
            .CK(us_clk), .Q(throttle_pwm_val_latched[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(123[14] 134[12])
    defparam throttle_pwm_val_latched__i4.GSR = "ENABLED";
    FD1P3AX throttle_pwm_val_latched__i5 (.D(\throttle_val[5] ), .SP(us_clk_enable_103), 
            .CK(us_clk), .Q(throttle_pwm_val_latched[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(123[14] 134[12])
    defparam throttle_pwm_val_latched__i5.GSR = "ENABLED";
    FD1P3AX throttle_pwm_val_latched__i6 (.D(\throttle_val[6] ), .SP(us_clk_enable_103), 
            .CK(us_clk), .Q(throttle_pwm_val_latched[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(123[14] 134[12])
    defparam throttle_pwm_val_latched__i6.GSR = "ENABLED";
    FD1P3AX throttle_pwm_val_latched__i7 (.D(\throttle_val[7] ), .SP(us_clk_enable_103), 
            .CK(us_clk), .Q(throttle_pwm_val_latched[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(123[14] 134[12])
    defparam throttle_pwm_val_latched__i7.GSR = "ENABLED";
    LUT4 i3_4_lut_adj_270 (.A(auto_state[2]), .B(auto_state[1]), .C(n52482), 
         .D(auto_state[3]), .Z(n44)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i3_4_lut_adj_270.init = 16'h0010;
    PFUMX i40906 (.BLUT(n52468), .ALUT(n52469), .C0(state[0]), .Z(next_state_4__N_1669));
    PFUMX i22769 (.BLUT(n48938), .ALUT(n48651), .C0(n8551), .Z(next_auto_state_8__N_1703));
    LUT4 i19912_3_lut (.A(n30583), .B(n30582), .C(n30524), .Z(count__auto_time_ms[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam i19912_3_lut.init = 16'hcaca;
    LUT4 i3_4_lut_adj_271 (.A(auto_state[4]), .B(n49305), .C(auto_state[5]), 
         .D(auto_state[3]), .Z(n8409)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (B+(C+!(D))))) */ ;
    defparam i3_4_lut_adj_271.init = 16'h0102;
    LUT4 i19921_3_lut_rep_490 (.A(n30592), .B(n30591), .C(n30524), .Z(n52426)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam i19921_3_lut_rep_490.init = 16'hcaca;
    LUT4 i1_2_lut_4_lut_adj_272 (.A(n30592), .B(n30591), .C(n30524), .D(count__auto_time_ms[27]), 
         .Z(n25)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam i1_2_lut_4_lut_adj_272.init = 16'hca00;
    LUT4 i23_1_lut (.A(state[3]), .Z(n17)) /* synthesis lut_function=(!(A)) */ ;
    defparam i23_1_lut.init = 16'h5555;
    LUT4 i7776_1_lut (.A(state[2]), .Z(n14)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(266[17:28])
    defparam i7776_1_lut.init = 16'h5555;
    LUT4 i29184_1_lut (.A(\next_state_4__N_1656[2] ), .Z(start_flag_N_1875)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(98[14] 105[42])
    defparam i29184_1_lut.init = 16'h5555;
    LUT4 i39840_4_lut (.A(n52213), .B(n4), .C(state[0]), .D(n48787), 
         .Z(n48533)) /* synthesis lut_function=(!((B (C+(D))+!B (C))+!A)) */ ;
    defparam i39840_4_lut.init = 16'h020a;
    LUT4 i16_4_lut (.A(state[2]), .B(n49347), .C(n52214), .D(n8_adj_5188), 
         .Z(n8)) /* synthesis lut_function=(!(A (B (C)+!B !((D)+!C))+!A (B+!(C (D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(154[17:51])
    defparam i16_4_lut.init = 16'h3a0a;
    LUT4 i38552_2_lut (.A(next_state[2]), .B(next_state[1]), .Z(n49347)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i38552_2_lut.init = 16'heeee;
    LUT4 i3_3_lut (.A(next_state[0]), .B(next_state[3]), .C(next_state[4]), 
         .Z(n8_adj_5188)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i3_3_lut.init = 16'h0404;
    LUT4 i1_2_lut_adj_273 (.A(us_clk_enable_66), .B(count__auto_time_ms_27__N_1767[27]), 
         .Z(n58[27])) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(69[15:34])
    defparam i1_2_lut_adj_273.init = 16'hdddd;
    LUT4 i2_3_lut_4_lut_adj_274 (.A(n52313), .B(n48170), .C(switch_b[0]), 
         .D(n52401), .Z(n48795)) /* synthesis lut_function=(!(A (C+!(D))+!A ((C+!(D))+!B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(159[53:84])
    defparam i2_3_lut_4_lut_adj_274.init = 16'h0e00;
    PFUMX mux_4101_i1 (.BLUT(n8620[0]), .ALUT(n48795), .C0(n8584), .Z(n8639[0]));
    LUT4 i1_2_lut_rep_253_3_lut_4_lut (.A(n52313), .B(n48170), .C(count__auto_time_ms[27]), 
         .D(\next_auto_state_8__N_1686[7] ), .Z(n52189)) /* synthesis lut_function=(A (C (D))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(159[53:84])
    defparam i1_2_lut_rep_253_3_lut_4_lut.init = 16'he000;
    LUT4 i37594_3_lut_4_lut (.A(state[2]), .B(state[1]), .C(state[3]), 
         .D(state[0]), .Z(n6)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;
    defparam i37594_3_lut_4_lut.init = 16'h0001;
    LUT4 i26944_2_lut_rep_499 (.A(state[3]), .B(state[2]), .Z(n52435)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i26944_2_lut_rep_499.init = 16'heeee;
    LUT4 i1_2_lut_rep_277_3_lut_4_lut (.A(state[3]), .B(state[2]), .C(state[4]), 
         .D(n52438), .Z(n52213)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i1_2_lut_rep_277_3_lut_4_lut.init = 16'h0100;
    LUT4 i1_4_lut_else_4_lut_adj_275 (.A(auto_state[5]), .B(auto_state[6]), 
         .C(auto_state[4]), .D(auto_state[7]), .Z(n52480)) /* synthesis lut_function=(!(A (B+(C+(D)))+!A (B (C+(D))+!B (C (D)+!C !(D))))) */ ;
    defparam i1_4_lut_else_4_lut_adj_275.init = 16'h0116;
    LUT4 i39644_3_lut (.A(state[4]), .B(n47358), .C(state[2]), .Z(next_state_4__N_1653)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(277[17:31])
    defparam i39644_3_lut.init = 16'h0202;
    LUT4 i2_3_lut_adj_276 (.A(state[0]), .B(state[3]), .C(state[1]), .Z(n47358)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(277[17:31])
    defparam i2_3_lut_adj_276.init = 16'hfefe;
    LUT4 i26890_2_lut (.A(state[4]), .B(state[1]), .Z(n37558)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i26890_2_lut.init = 16'heeee;
    LUT4 count__auto_time_ms_i1_i27_3_lut (.A(count__auto_time_ms[26]), .B(count__auto_time_ms_27__N_1767[26]), 
         .C(us_clk_enable_66), .Z(n58[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i1_i27_3_lut.init = 16'hcaca;
    LUT4 i19858_3_lut (.A(n30529), .B(n30528), .C(n30524), .Z(count__auto_time_ms[26])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam i19858_3_lut.init = 16'hcaca;
    LUT4 i39850_4_lut (.A(n45_adj_5189), .B(n37_adj_5190), .C(n44_adj_5191), 
         .D(n38_adj_5192), .Z(us_clk_enable_66)) /* synthesis lut_function=(!(A (B (C (D))))) */ ;
    defparam i39850_4_lut.init = 16'h7fff;
    LUT4 i21_4_lut (.A(count__auto_time_ms[16]), .B(n42_adj_5193), .C(n34), 
         .D(count__auto_time_ms[20]), .Z(n45_adj_5189)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i21_4_lut.init = 16'h8000;
    LUT4 i13_4_lut (.A(n25), .B(n7_adj_5194), .C(count__auto_time_ms[6]), 
         .D(n8_adj_5195), .Z(n37_adj_5190)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i13_4_lut.init = 16'h8000;
    LUT4 i20_4_lut (.A(count__auto_time_ms[3]), .B(n40_adj_5196), .C(n30), 
         .D(count__auto_time_ms[11]), .Z(n44_adj_5191)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i20_4_lut.init = 16'h8000;
    LUT4 i14_4_lut (.A(count__auto_time_ms[15]), .B(count__auto_time_ms[18]), 
         .C(count__auto_time_ms[24]), .D(count__auto_time_ms[17]), .Z(n38_adj_5192)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i14_4_lut.init = 16'h8000;
    LUT4 i18_4_lut (.A(count__auto_time_ms[12]), .B(count__auto_time_ms[5]), 
         .C(count__auto_time_ms[23]), .D(count__auto_time_ms[26]), .Z(n42_adj_5193)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i18_4_lut.init = 16'h8000;
    LUT4 i2_2_lut (.A(count__auto_time_ms[10]), .B(count__auto_time_ms[8]), 
         .Z(n7_adj_5194)) /* synthesis lut_function=(A (B)) */ ;
    defparam i2_2_lut.init = 16'h8888;
    LUT4 i3_3_lut_adj_277 (.A(count__auto_time_ms[13]), .B(count__auto_time_ms[4]), 
         .C(count__auto_time_ms[9]), .Z(n8_adj_5195)) /* synthesis lut_function=(A (B (C))) */ ;
    defparam i3_3_lut_adj_277.init = 16'h8080;
    LUT4 i16_4_lut_adj_278 (.A(count__auto_time_ms[22]), .B(count__auto_time_ms[14]), 
         .C(count__auto_time_ms[21]), .D(count__auto_time_ms[1]), .Z(n40_adj_5196)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i16_4_lut_adj_278.init = 16'h8000;
    LUT4 i19870_3_lut (.A(n30541), .B(n30540), .C(n30524), .Z(count__auto_time_ms[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam i19870_3_lut.init = 16'hcaca;
    LUT4 i19894_3_lut (.A(n30565), .B(n30564), .C(n30524), .Z(count__auto_time_ms[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam i19894_3_lut.init = 16'hcaca;
    LUT4 i19873_3_lut (.A(n30544), .B(n30543), .C(n30524), .Z(count__auto_time_ms[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam i19873_3_lut.init = 16'hcaca;
    LUT4 i19903_3_lut (.A(n30574), .B(n30573), .C(n30524), .Z(count__auto_time_ms[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam i19903_3_lut.init = 16'hcaca;
    LUT4 i19897_3_lut (.A(n30568), .B(n30567), .C(n30524), .Z(count__auto_time_ms[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam i19897_3_lut.init = 16'hcaca;
    LUT4 i19909_3_lut (.A(n30580), .B(n30579), .C(n30524), .Z(count__auto_time_ms[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam i19909_3_lut.init = 16'hcaca;
    LUT4 i19867_3_lut (.A(n30538), .B(n30537), .C(n30524), .Z(count__auto_time_ms[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam i19867_3_lut.init = 16'hcaca;
    LUT4 i19891_3_lut (.A(n30562), .B(n30561), .C(n30524), .Z(count__auto_time_ms[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam i19891_3_lut.init = 16'hcaca;
    LUT4 i19882_3_lut (.A(n30553), .B(n30552), .C(n30524), .Z(count__auto_time_ms[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam i19882_3_lut.init = 16'hcaca;
    LUT4 i19864_3_lut (.A(n30535), .B(n30534), .C(n30524), .Z(count__auto_time_ms[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam i19864_3_lut.init = 16'hcaca;
    LUT4 i19885_3_lut (.A(n30556), .B(n30555), .C(n30524), .Z(count__auto_time_ms[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam i19885_3_lut.init = 16'hcaca;
    LUT4 i19900_3_lut (.A(n30571), .B(n30570), .C(n30524), .Z(count__auto_time_ms[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam i19900_3_lut.init = 16'hcaca;
    LUT4 i19906_3_lut (.A(n30577), .B(n30576), .C(n30524), .Z(count__auto_time_ms[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam i19906_3_lut.init = 16'hcaca;
    LUT4 i19888_3_lut (.A(n30559), .B(n30558), .C(n30524), .Z(count__auto_time_ms[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam i19888_3_lut.init = 16'hcaca;
    LUT4 i19876_3_lut (.A(n30547), .B(n30546), .C(n30524), .Z(count__auto_time_ms[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam i19876_3_lut.init = 16'hcaca;
    LUT4 count__auto_time_ms_i1_i26_3_lut (.A(n52326), .B(count__auto_time_ms_27__N_1767[25]), 
         .C(us_clk_enable_66), .Z(n58[25])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i1_i26_3_lut.init = 16'hcaca;
    LUT4 count__auto_time_ms_i1_i25_3_lut (.A(count__auto_time_ms[24]), .B(count__auto_time_ms_27__N_1767[24]), 
         .C(us_clk_enable_66), .Z(n58[24])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i1_i25_3_lut.init = 16'hcaca;
    LUT4 count__auto_time_ms_i1_i24_3_lut (.A(count__auto_time_ms[23]), .B(count__auto_time_ms_27__N_1767[23]), 
         .C(us_clk_enable_66), .Z(n58[23])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i1_i24_3_lut.init = 16'hcaca;
    LUT4 count__auto_time_ms_i1_i23_3_lut (.A(count__auto_time_ms[22]), .B(count__auto_time_ms_27__N_1767[22]), 
         .C(us_clk_enable_66), .Z(n58[22])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i1_i23_3_lut.init = 16'hcaca;
    LUT4 count__auto_time_ms_i1_i22_3_lut (.A(count__auto_time_ms[21]), .B(count__auto_time_ms_27__N_1767[21]), 
         .C(us_clk_enable_66), .Z(n58[21])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i1_i22_3_lut.init = 16'hcaca;
    LUT4 count__auto_time_ms_i1_i21_3_lut (.A(count__auto_time_ms[20]), .B(count__auto_time_ms_27__N_1767[20]), 
         .C(us_clk_enable_66), .Z(n58[20])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i1_i21_3_lut.init = 16'hcaca;
    LUT4 count__auto_time_ms_i1_i20_3_lut (.A(n52325), .B(count__auto_time_ms_27__N_1767[19]), 
         .C(us_clk_enable_66), .Z(n58[19])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i1_i20_3_lut.init = 16'hcaca;
    LUT4 count__auto_time_ms_i1_i19_3_lut (.A(count__auto_time_ms[18]), .B(count__auto_time_ms_27__N_1767[18]), 
         .C(us_clk_enable_66), .Z(n58[18])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i1_i19_3_lut.init = 16'hcaca;
    LUT4 count__auto_time_ms_i1_i18_3_lut (.A(count__auto_time_ms[17]), .B(count__auto_time_ms_27__N_1767[17]), 
         .C(us_clk_enable_66), .Z(n58[17])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i1_i18_3_lut.init = 16'hcaca;
    LUT4 count__auto_time_ms_i1_i17_3_lut (.A(count__auto_time_ms[16]), .B(count__auto_time_ms_27__N_1767[16]), 
         .C(us_clk_enable_66), .Z(n58[16])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i1_i17_3_lut.init = 16'hcaca;
    LUT4 count__auto_time_ms_i1_i16_3_lut (.A(count__auto_time_ms[15]), .B(count__auto_time_ms_27__N_1767[15]), 
         .C(us_clk_enable_66), .Z(n58[15])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i1_i16_3_lut.init = 16'hcaca;
    LUT4 count__auto_time_ms_i1_i15_3_lut (.A(count__auto_time_ms[14]), .B(count__auto_time_ms_27__N_1767[14]), 
         .C(us_clk_enable_66), .Z(n58[14])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i1_i15_3_lut.init = 16'hcaca;
    LUT4 count__auto_time_ms_i1_i13_3_lut (.A(count__auto_time_ms[12]), .B(count__auto_time_ms_27__N_1767[12]), 
         .C(us_clk_enable_66), .Z(n58[12])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i1_i13_3_lut.init = 16'hcaca;
    LUT4 count__auto_time_ms_i1_i12_3_lut (.A(count__auto_time_ms[11]), .B(count__auto_time_ms_27__N_1767[11]), 
         .C(us_clk_enable_66), .Z(n58[11])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i1_i12_3_lut.init = 16'hcaca;
    LUT4 count__auto_time_ms_i1_i8_3_lut (.A(count__auto_time_ms[7]), .B(count__auto_time_ms_27__N_1767[7]), 
         .C(us_clk_enable_66), .Z(n58[7])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i1_i8_3_lut.init = 16'hcaca;
    LUT4 count__auto_time_ms_i1_i7_3_lut (.A(count__auto_time_ms[6]), .B(count__auto_time_ms_27__N_1767[6]), 
         .C(us_clk_enable_66), .Z(n58[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i1_i7_3_lut.init = 16'hcaca;
    LUT4 count__auto_time_ms_i1_i6_3_lut (.A(count__auto_time_ms[5]), .B(count__auto_time_ms_27__N_1767[5]), 
         .C(us_clk_enable_66), .Z(n58[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i1_i6_3_lut.init = 16'hcaca;
    LUT4 count__auto_time_ms_i1_i4_3_lut (.A(count__auto_time_ms[3]), .B(count__auto_time_ms_27__N_1767[3]), 
         .C(us_clk_enable_66), .Z(n58[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i1_i4_3_lut.init = 16'hcaca;
    LUT4 count__auto_time_ms_i1_i3_3_lut (.A(count__auto_time_ms[2]), .B(count__auto_time_ms_27__N_1767[2]), 
         .C(us_clk_enable_66), .Z(n58[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i1_i3_3_lut.init = 16'hcaca;
    LUT4 count__auto_time_ms_i1_i2_3_lut (.A(count__auto_time_ms[1]), .B(count__auto_time_ms_27__N_1767[1]), 
         .C(us_clk_enable_66), .Z(n58[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i1_i2_3_lut.init = 16'hcaca;
    LUT4 count__auto_time_ms_i1_i1_3_lut (.A(n52426), .B(count__auto_time_ms_27__N_1767[0]), 
         .C(us_clk_enable_66), .Z(n58[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i1_i1_3_lut.init = 16'hcaca;
    CCU2D sub_8_add_2_29 (.A0(count__auto_time_ms[27]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n43834), .S0(count__auto_time_ms_27__N_1767[27]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(90[36:64])
    defparam sub_8_add_2_29.INIT0 = 16'h5555;
    defparam sub_8_add_2_29.INIT1 = 16'h0000;
    defparam sub_8_add_2_29.INJECT1_0 = "NO";
    defparam sub_8_add_2_29.INJECT1_1 = "NO";
    CCU2D sub_8_add_2_27 (.A0(n52326), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count__auto_time_ms[26]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n43833), .COUT(n43834), .S0(count__auto_time_ms_27__N_1767[25]), 
          .S1(count__auto_time_ms_27__N_1767[26]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(90[36:64])
    defparam sub_8_add_2_27.INIT0 = 16'h5555;
    defparam sub_8_add_2_27.INIT1 = 16'h5555;
    defparam sub_8_add_2_27.INJECT1_0 = "NO";
    defparam sub_8_add_2_27.INJECT1_1 = "NO";
    CCU2D sub_8_add_2_25 (.A0(count__auto_time_ms[23]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count__auto_time_ms[24]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43832), .COUT(n43833), .S0(count__auto_time_ms_27__N_1767[23]), 
          .S1(count__auto_time_ms_27__N_1767[24]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(90[36:64])
    defparam sub_8_add_2_25.INIT0 = 16'h5555;
    defparam sub_8_add_2_25.INIT1 = 16'h5555;
    defparam sub_8_add_2_25.INJECT1_0 = "NO";
    defparam sub_8_add_2_25.INJECT1_1 = "NO";
    CCU2D sub_8_add_2_23 (.A0(count__auto_time_ms[21]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count__auto_time_ms[22]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43831), .COUT(n43832), .S0(count__auto_time_ms_27__N_1767[21]), 
          .S1(count__auto_time_ms_27__N_1767[22]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(90[36:64])
    defparam sub_8_add_2_23.INIT0 = 16'h5555;
    defparam sub_8_add_2_23.INIT1 = 16'h5555;
    defparam sub_8_add_2_23.INJECT1_0 = "NO";
    defparam sub_8_add_2_23.INJECT1_1 = "NO";
    LUT4 i12_4_lut (.A(n19), .B(n24), .C(next_state[2]), .D(n14_adj_5197), 
         .Z(n33315)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(138[5] 228[8])
    defparam i12_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(next_state[4]), .B(auto_state[1]), .Z(n19)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(138[5] 228[8])
    defparam i6_2_lut.init = 16'heeee;
    LUT4 i11_4_lut (.A(next_state[0]), .B(n22), .C(n16), .D(auto_state[6]), 
         .Z(n24)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(138[5] 228[8])
    defparam i11_4_lut.init = 16'hfffe;
    LUT4 i22777_3_lut_4_lut_4_lut (.A(n52237), .B(\next_auto_state_8__N_1686[7] ), 
         .C(auto_state[0]), .D(count__auto_time_ms[27]), .Z(n8620[0])) /* synthesis lut_function=(A (B (C+(D))+!B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(123[14] 134[12])
    defparam i22777_3_lut_4_lut_4_lut.init = 16'ha8a0;
    LUT4 i1_3_lut (.A(auto_state[5]), .B(auto_state[3]), .C(auto_state[4]), 
         .Z(n14_adj_5197)) /* synthesis lut_function=(A+(B (C)+!B !(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(138[5] 228[8])
    defparam i1_3_lut.init = 16'hebeb;
    CCU2D sub_8_add_2_21 (.A0(n52325), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(count__auto_time_ms[20]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n43830), .COUT(n43831), .S0(count__auto_time_ms_27__N_1767[19]), 
          .S1(count__auto_time_ms_27__N_1767[20]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(90[36:64])
    defparam sub_8_add_2_21.INIT0 = 16'h5555;
    defparam sub_8_add_2_21.INIT1 = 16'h5555;
    defparam sub_8_add_2_21.INJECT1_0 = "NO";
    defparam sub_8_add_2_21.INJECT1_1 = "NO";
    LUT4 i9_4_lut (.A(next_state[1]), .B(next_state[3]), .C(auto_state[8]), 
         .D(auto_state[7]), .Z(n22)) /* synthesis lut_function=(A+((C+(D))+!B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(138[5] 228[8])
    defparam i9_4_lut.init = 16'hfffb;
    LUT4 i3_2_lut (.A(auto_state[2]), .B(auto_state[0]), .Z(n16)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(138[5] 228[8])
    defparam i3_2_lut.init = 16'heeee;
    PFUMX i40974 (.BLUT(n52570), .ALUT(n52571), .C0(state[0]), .Z(n52572));
    CCU2D sub_8_add_2_19 (.A0(count__auto_time_ms[17]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count__auto_time_ms[18]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43829), .COUT(n43830), .S0(count__auto_time_ms_27__N_1767[17]), 
          .S1(count__auto_time_ms_27__N_1767[18]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(90[36:64])
    defparam sub_8_add_2_19.INIT0 = 16'h5555;
    defparam sub_8_add_2_19.INIT1 = 16'h5555;
    defparam sub_8_add_2_19.INJECT1_0 = "NO";
    defparam sub_8_add_2_19.INJECT1_1 = "NO";
    PFUMX i40543 (.BLUT(n51604), .ALUT(n51603), .C0(n8551), .Z(n51605));
    CCU2D sub_8_add_2_17 (.A0(count__auto_time_ms[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count__auto_time_ms[16]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43828), .COUT(n43829), .S0(count__auto_time_ms_27__N_1767[15]), 
          .S1(count__auto_time_ms_27__N_1767[16]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(90[36:64])
    defparam sub_8_add_2_17.INIT0 = 16'h5555;
    defparam sub_8_add_2_17.INIT1 = 16'h5555;
    defparam sub_8_add_2_17.INJECT1_0 = "NO";
    defparam sub_8_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_8_add_2_15 (.A0(count__auto_time_ms[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count__auto_time_ms[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43827), .COUT(n43828), .S0(count__auto_time_ms_27__N_1767[13]), 
          .S1(count__auto_time_ms_27__N_1767[14]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(90[36:64])
    defparam sub_8_add_2_15.INIT0 = 16'h5555;
    defparam sub_8_add_2_15.INIT1 = 16'h5555;
    defparam sub_8_add_2_15.INJECT1_0 = "NO";
    defparam sub_8_add_2_15.INJECT1_1 = "NO";
    CCU2D sub_8_add_2_13 (.A0(count__auto_time_ms[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count__auto_time_ms[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43826), .COUT(n43827), .S0(count__auto_time_ms_27__N_1767[11]), 
          .S1(count__auto_time_ms_27__N_1767[12]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(90[36:64])
    defparam sub_8_add_2_13.INIT0 = 16'h5555;
    defparam sub_8_add_2_13.INIT1 = 16'h5555;
    defparam sub_8_add_2_13.INJECT1_0 = "NO";
    defparam sub_8_add_2_13.INJECT1_1 = "NO";
    CCU2D sub_8_add_2_11 (.A0(count__auto_time_ms[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count__auto_time_ms[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43825), .COUT(n43826), .S0(count__auto_time_ms_27__N_1767[9]), 
          .S1(count__auto_time_ms_27__N_1767[10]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(90[36:64])
    defparam sub_8_add_2_11.INIT0 = 16'h5555;
    defparam sub_8_add_2_11.INIT1 = 16'h5555;
    defparam sub_8_add_2_11.INJECT1_0 = "NO";
    defparam sub_8_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_8_add_2_9 (.A0(count__auto_time_ms[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count__auto_time_ms[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43824), .COUT(n43825), .S0(count__auto_time_ms_27__N_1767[7]), 
          .S1(count__auto_time_ms_27__N_1767[8]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(90[36:64])
    defparam sub_8_add_2_9.INIT0 = 16'h5555;
    defparam sub_8_add_2_9.INIT1 = 16'h5555;
    defparam sub_8_add_2_9.INJECT1_0 = "NO";
    defparam sub_8_add_2_9.INJECT1_1 = "NO";
    FD1S1I next_state_4__I_50_i5 (.D(n52566), .CK(next_state_4__N_1669), 
           .CD(n17), .Q(next_state[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(138[5] 228[8])
    defparam next_state_4__I_50_i5.GSR = "ENABLED";
    FD1S1I next_state_4__I_50_i4 (.D(n51), .CK(next_state_4__N_1669), .CD(n14), 
           .Q(next_state[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(138[5] 228[8])
    defparam next_state_4__I_50_i4.GSR = "ENABLED";
    FD1S1I next_state_4__I_50_i3 (.D(n48533), .CK(next_state_4__N_1669), 
           .CD(start_flag_N_1875), .Q(next_state[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(138[5] 228[8])
    defparam next_state_4__I_50_i3.GSR = "ENABLED";
    FD1S3DX count__auto_time_ms_i0_i0_19919_19920_reset (.D(n58[0]), .CK(us_clk), 
            .CD(count__auto_time_ms_27__N_1647), .Q(n30592)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i0_19919_19920_reset.GSR = "DISABLED";
    FD1S3DX count__auto_time_ms_i0_i1_19916_19917_reset (.D(n58[1]), .CK(us_clk), 
            .CD(count__auto_time_ms_27__N_1647), .Q(n30589)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i1_19916_19917_reset.GSR = "DISABLED";
    FD1S3DX count__auto_time_ms_i0_i2_19913_19914_reset (.D(n58[2]), .CK(us_clk), 
            .CD(count__auto_time_ms_27__N_1647), .Q(n30586)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i2_19913_19914_reset.GSR = "DISABLED";
    FD1S3DX count__auto_time_ms_i0_i3_19910_19911_reset (.D(n58[3]), .CK(us_clk), 
            .CD(count__auto_time_ms_27__N_1647), .Q(n30583)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i3_19910_19911_reset.GSR = "DISABLED";
    FD1S3DX count__auto_time_ms_i0_i5_19907_19908_reset (.D(n58[5]), .CK(us_clk), 
            .CD(count__auto_time_ms_27__N_1647), .Q(n30580)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i5_19907_19908_reset.GSR = "DISABLED";
    FD1S3DX count__auto_time_ms_i0_i6_19904_19905_reset (.D(n58[6]), .CK(us_clk), 
            .CD(count__auto_time_ms_27__N_1647), .Q(n30577)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i6_19904_19905_reset.GSR = "DISABLED";
    FD1S3DX count__auto_time_ms_i0_i7_19901_19902_reset (.D(n58[7]), .CK(us_clk), 
            .CD(count__auto_time_ms_27__N_1647), .Q(n30574)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i7_19901_19902_reset.GSR = "DISABLED";
    FD1S3DX count__auto_time_ms_i0_i11_19898_19899_reset (.D(n58[11]), .CK(us_clk), 
            .CD(count__auto_time_ms_27__N_1647), .Q(n30571)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i11_19898_19899_reset.GSR = "DISABLED";
    FD1S3DX count__auto_time_ms_i0_i12_19895_19896_reset (.D(n58[12]), .CK(us_clk), 
            .CD(count__auto_time_ms_27__N_1647), .Q(n30568)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i12_19895_19896_reset.GSR = "DISABLED";
    FD1S3DX count__auto_time_ms_i0_i14_19892_19893_reset (.D(n58[14]), .CK(us_clk), 
            .CD(count__auto_time_ms_27__N_1647), .Q(n30565)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i14_19892_19893_reset.GSR = "DISABLED";
    FD1S3DX count__auto_time_ms_i0_i15_19889_19890_reset (.D(n58[15]), .CK(us_clk), 
            .CD(count__auto_time_ms_27__N_1647), .Q(n30562)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i15_19889_19890_reset.GSR = "DISABLED";
    FD1S3DX count__auto_time_ms_i0_i16_19886_19887_reset (.D(n58[16]), .CK(us_clk), 
            .CD(count__auto_time_ms_27__N_1647), .Q(n30559)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i16_19886_19887_reset.GSR = "DISABLED";
    FD1S3DX count__auto_time_ms_i0_i17_19883_19884_reset (.D(n58[17]), .CK(us_clk), 
            .CD(count__auto_time_ms_27__N_1647), .Q(n30556)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i17_19883_19884_reset.GSR = "DISABLED";
    FD1S3DX count__auto_time_ms_i0_i18_19880_19881_reset (.D(n58[18]), .CK(us_clk), 
            .CD(count__auto_time_ms_27__N_1647), .Q(n30553)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i18_19880_19881_reset.GSR = "DISABLED";
    FD1S3DX count__auto_time_ms_i0_i19_19877_19878_reset (.D(n58[19]), .CK(us_clk), 
            .CD(count__auto_time_ms_27__N_1647), .Q(n30550)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i19_19877_19878_reset.GSR = "DISABLED";
    FD1S3DX count__auto_time_ms_i0_i20_19874_19875_reset (.D(n58[20]), .CK(us_clk), 
            .CD(count__auto_time_ms_27__N_1647), .Q(n30547)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i20_19874_19875_reset.GSR = "DISABLED";
    FD1S3DX count__auto_time_ms_i0_i21_19871_19872_reset (.D(n58[21]), .CK(us_clk), 
            .CD(count__auto_time_ms_27__N_1647), .Q(n30544)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i21_19871_19872_reset.GSR = "DISABLED";
    FD1S3DX count__auto_time_ms_i0_i22_19868_19869_reset (.D(n58[22]), .CK(us_clk), 
            .CD(count__auto_time_ms_27__N_1647), .Q(n30541)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i22_19868_19869_reset.GSR = "DISABLED";
    FD1S3DX count__auto_time_ms_i0_i23_19865_19866_reset (.D(n58[23]), .CK(us_clk), 
            .CD(count__auto_time_ms_27__N_1647), .Q(n30538)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i23_19865_19866_reset.GSR = "DISABLED";
    FD1S3DX count__auto_time_ms_i0_i24_19862_19863_reset (.D(n58[24]), .CK(us_clk), 
            .CD(count__auto_time_ms_27__N_1647), .Q(n30535)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i24_19862_19863_reset.GSR = "DISABLED";
    FD1S3DX count__auto_time_ms_i0_i25_19859_19860_reset (.D(n58[25]), .CK(us_clk), 
            .CD(count__auto_time_ms_27__N_1647), .Q(n30532)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i25_19859_19860_reset.GSR = "DISABLED";
    FD1S3DX count__auto_time_ms_i0_i26_19856_19857_reset (.D(n58[26]), .CK(us_clk), 
            .CD(count__auto_time_ms_27__N_1647), .Q(n30529)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i26_19856_19857_reset.GSR = "DISABLED";
    FD1S3DX count__auto_time_ms_i0_i27_19853_19854_reset (.D(n58[27]), .CK(us_clk), 
            .CD(count__auto_time_ms_27__N_1647), .Q(n30526)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i27_19853_19854_reset.GSR = "DISABLED";
    FD1S3AY count__auto_time_ms_i0_i27_19853_19854_set (.D(n58[27]), .CK(us_clk), 
            .Q(n30525)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=26, LSE_RCOL=6, LSE_LLINE=362, LSE_RLINE=375 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(89[14] 90[65])
    defparam count__auto_time_ms_i0_i27_19853_19854_set.GSR = "ENABLED";
    CCU2D sub_8_add_2_7 (.A0(count__auto_time_ms[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(count__auto_time_ms[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43823), .COUT(n43824), .S0(count__auto_time_ms_27__N_1767[5]), 
          .S1(count__auto_time_ms_27__N_1767[6]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/auto_mode_controller.v(90[36:64])
    defparam sub_8_add_2_7.INIT0 = 16'h5555;
    defparam sub_8_add_2_7.INIT1 = 16'h5555;
    defparam sub_8_add_2_7.INJECT1_0 = "NO";
    defparam sub_8_add_2_7.INJECT1_1 = "NO";
    
endmodule
//
// Verilog Description of module flight_mode
//

module flight_mode (switch_b, us_clk, \swa_swb_val[7] , \swa_swb_val[4] , 
            \swa_swb_val[5] , \swa_swb_val[3] , \swa_swb_val[6] , \swa_swb_val[2] , 
            n10, \next_auto_state_8__N_1686[7] , n52359, \swa_swb_val[1] ) /* synthesis syn_module_defined=1 */ ;
    output [1:0]switch_b;
    input us_clk;
    input \swa_swb_val[7] ;
    input \swa_swb_val[4] ;
    input \swa_swb_val[5] ;
    input \swa_swb_val[3] ;
    input \swa_swb_val[6] ;
    input \swa_swb_val[2] ;
    input n10;
    output \next_auto_state_8__N_1686[7] ;
    input n52359;
    input \swa_swb_val[1] ;
    
    wire us_clk /* synthesis SET_AS_NETWORK=us_clk, is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(221[10:16])
    wire [1:0]switch_b_1__N_274;
    
    wire n48464, n38173, n52055, switch_a_2__N_283, switch_a_2__N_279, 
        n10_c, n7, n4, n50402, n48659;
    wire [2:0]switch_a_2__N_269;
    
    wire n6, n6_adj_5178;
    
    FD1S3AX switch_b_i0 (.D(switch_b_1__N_274[0]), .CK(us_clk), .Q(switch_b[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=287 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/flight_mode.v(30[14] 39[12])
    defparam switch_b_i0.GSR = "ENABLED";
    LUT4 i37678_4_lut (.A(\swa_swb_val[7] ), .B(\swa_swb_val[4] ), .C(\swa_swb_val[5] ), 
         .D(\swa_swb_val[3] ), .Z(n48464)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i37678_4_lut.init = 16'haaa8;
    LUT4 n38173_bdd_3_lut (.A(n38173), .B(\swa_swb_val[7] ), .C(\swa_swb_val[6] ), 
         .Z(n52055)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam n38173_bdd_3_lut.init = 16'h2020;
    LUT4 i2_4_lut (.A(switch_a_2__N_283), .B(switch_a_2__N_279), .C(\swa_swb_val[7] ), 
         .D(n10_c), .Z(switch_b_1__N_274[0])) /* synthesis lut_function=(A+!(B ((D)+!C))) */ ;
    defparam i2_4_lut.init = 16'hbbfb;
    LUT4 i4_4_lut (.A(n7), .B(n48464), .C(\swa_swb_val[5] ), .D(n4), 
         .Z(n10_c)) /* synthesis lut_function=(A+!(B (C+(D)))) */ ;
    defparam i4_4_lut.init = 16'hbbbf;
    LUT4 i1_4_lut (.A(\swa_swb_val[6] ), .B(n50402), .C(n48659), .D(\swa_swb_val[5] ), 
         .Z(n7)) /* synthesis lut_function=((B (C (D))+!B (C+!(D)))+!A) */ ;
    defparam i1_4_lut.init = 16'hf577;
    LUT4 n4_bdd_4_lut (.A(n4), .B(\swa_swb_val[7] ), .C(n52055), .D(\swa_swb_val[5] ), 
         .Z(switch_a_2__N_283)) /* synthesis lut_function=(A (C (D))+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam n4_bdd_4_lut.init = 16'hf044;
    LUT4 i1_rep_8_2_lut (.A(\swa_swb_val[3] ), .B(\swa_swb_val[4] ), .Z(n50402)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_rep_8_2_lut.init = 16'heeee;
    LUT4 i2_4_lut_adj_252 (.A(\swa_swb_val[4] ), .B(\swa_swb_val[2] ), .C(\swa_swb_val[3] ), 
         .D(n10), .Z(n48659)) /* synthesis lut_function=(A (B (C)+!B (C (D)))) */ ;
    defparam i2_4_lut_adj_252.init = 16'ha080;
    FD1S3AX switch_a_i2 (.D(switch_a_2__N_269[2]), .CK(us_clk), .Q(\next_auto_state_8__N_1686[7] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=287 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/flight_mode.v(30[14] 39[12])
    defparam switch_a_i2.GSR = "ENABLED";
    FD1S3AX switch_b_i1 (.D(switch_b_1__N_274[1]), .CK(us_clk), .Q(switch_b[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=17, LSE_RCOL=6, LSE_LLINE=281, LSE_RLINE=287 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/flight_mode.v(30[14] 39[12])
    defparam switch_b_i1.GSR = "ENABLED";
    LUT4 i2_3_lut (.A(n6), .B(\swa_swb_val[7] ), .C(\swa_swb_val[6] ), 
         .Z(switch_a_2__N_279)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut.init = 16'hfefe;
    LUT4 i2_4_lut_adj_253 (.A(\swa_swb_val[4] ), .B(\swa_swb_val[5] ), .C(\swa_swb_val[3] ), 
         .D(n52359), .Z(n6)) /* synthesis lut_function=(A (B (C+(D)))) */ ;
    defparam i2_4_lut_adj_253.init = 16'h8880;
    LUT4 i1_4_lut_adj_254 (.A(\swa_swb_val[6] ), .B(n6_adj_5178), .C(\swa_swb_val[4] ), 
         .D(\swa_swb_val[3] ), .Z(n4)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;
    defparam i1_4_lut_adj_254.init = 16'hfaea;
    LUT4 i7174_2_lut (.A(\swa_swb_val[1] ), .B(\swa_swb_val[2] ), .Z(n6_adj_5178)) /* synthesis lut_function=(A (B)) */ ;
    defparam i7174_2_lut.init = 16'h8888;
    LUT4 i39768_4_lut (.A(\swa_swb_val[7] ), .B(n38173), .C(\swa_swb_val[6] ), 
         .D(\swa_swb_val[5] ), .Z(switch_a_2__N_269[2])) /* synthesis lut_function=(!(A+(B (C (D))))) */ ;
    defparam i39768_4_lut.init = 16'h1555;
    LUT4 i27473_3_lut (.A(\swa_swb_val[2] ), .B(\swa_swb_val[3] ), .C(\swa_swb_val[4] ), 
         .Z(n38173)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i27473_3_lut.init = 16'hfefe;
    LUT4 i25_4_lut (.A(\swa_swb_val[7] ), .B(n48464), .C(\swa_swb_val[6] ), 
         .D(n6), .Z(switch_b_1__N_274[1])) /* synthesis lut_function=(!(A (B (C))+!A (B (C+!(D))+!B !(C+(D))))) */ ;
    defparam i25_4_lut.init = 16'h3f3a;
    
endmodule
//
// Verilog Description of module pwm_generator
//

module pwm_generator (us_clk, us_clk_enable_61, high_counter_9__N_4408, 
            \next_state_2__N_4443[0] , GND_net, n53885, resetn, motor_4_pwm_c, 
            motor_3_pwm_c, motor_2_pwm_c, motor_1_pwm_c) /* synthesis syn_module_defined=1 */ ;
    input us_clk;
    input us_clk_enable_61;
    output high_counter_9__N_4408;
    output \next_state_2__N_4443[0] ;
    input GND_net;
    input n53885;
    input resetn;
    output motor_4_pwm_c;
    output motor_3_pwm_c;
    output motor_2_pwm_c;
    output motor_1_pwm_c;
    
    wire us_clk /* synthesis SET_AS_NETWORK=us_clk, is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(221[10:16])
    wire [9:0]high_counter;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(48[39:51])
    wire [9:0]n29;
    wire [15:0]period_counter;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(47[16:30])
    wire [15:0]period_counter_15__N_4409;
    
    wire n30656;
    wire [15:0]n1;
    
    wire n43819, n43818, n43817, n43816, high_counter_en, n27989, 
        n8, n14_adj_5175, n10, n52406, n11, n9, n43814, n7, 
        n7_adj_5176, n47352, n52405, n43813, n43812, n43811, n43810, 
        n43809, n43808, n43807;
    wire [2:0]next_state_2__N_4440;
    
    wire n48020, n36457, n48749;
    
    FD1P3IX high_counter__i0 (.D(n29[0]), .SP(us_clk_enable_61), .CD(high_counter_9__N_4408), 
            .CK(us_clk), .Q(high_counter[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=19, LSE_RCOL=25, LSE_LLINE=495, LSE_RLINE=507 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(112[14] 131[12])
    defparam high_counter__i0.GSR = "ENABLED";
    FD1S3IX period_counter__i0 (.D(period_counter_15__N_4409[0]), .CK(us_clk), 
            .CD(high_counter_9__N_4408), .Q(period_counter[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=19, LSE_RCOL=25, LSE_LLINE=495, LSE_RLINE=507 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(112[14] 131[12])
    defparam period_counter__i0.GSR = "ENABLED";
    FD1S3IX period_counter__i14 (.D(n1[14]), .CK(us_clk), .CD(n30656), 
            .Q(period_counter[14])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=19, LSE_RCOL=25, LSE_LLINE=495, LSE_RLINE=507 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(112[14] 131[12])
    defparam period_counter__i14.GSR = "ENABLED";
    FD1S3IX period_counter__i13 (.D(n1[13]), .CK(us_clk), .CD(n30656), 
            .Q(period_counter[13])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=19, LSE_RCOL=25, LSE_LLINE=495, LSE_RLINE=507 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(112[14] 131[12])
    defparam period_counter__i13.GSR = "ENABLED";
    FD1S3IX period_counter__i12 (.D(n1[12]), .CK(us_clk), .CD(n30656), 
            .Q(period_counter[12])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=19, LSE_RCOL=25, LSE_LLINE=495, LSE_RLINE=507 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(112[14] 131[12])
    defparam period_counter__i12.GSR = "ENABLED";
    FD1S3IX period_counter__i11 (.D(n1[11]), .CK(us_clk), .CD(n30656), 
            .Q(period_counter[11])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=19, LSE_RCOL=25, LSE_LLINE=495, LSE_RLINE=507 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(112[14] 131[12])
    defparam period_counter__i11.GSR = "ENABLED";
    FD1S3IX period_counter__i10 (.D(n1[10]), .CK(us_clk), .CD(n30656), 
            .Q(period_counter[10])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=19, LSE_RCOL=25, LSE_LLINE=495, LSE_RLINE=507 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(112[14] 131[12])
    defparam period_counter__i10.GSR = "ENABLED";
    FD1S3IX period_counter__i9 (.D(period_counter_15__N_4409[9]), .CK(us_clk), 
            .CD(high_counter_9__N_4408), .Q(period_counter[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=19, LSE_RCOL=25, LSE_LLINE=495, LSE_RLINE=507 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(112[14] 131[12])
    defparam period_counter__i9.GSR = "ENABLED";
    FD1S3IX period_counter__i8 (.D(period_counter_15__N_4409[8]), .CK(us_clk), 
            .CD(high_counter_9__N_4408), .Q(period_counter[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=19, LSE_RCOL=25, LSE_LLINE=495, LSE_RLINE=507 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(112[14] 131[12])
    defparam period_counter__i8.GSR = "ENABLED";
    FD1S3IX period_counter__i7 (.D(period_counter_15__N_4409[7]), .CK(us_clk), 
            .CD(high_counter_9__N_4408), .Q(period_counter[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=19, LSE_RCOL=25, LSE_LLINE=495, LSE_RLINE=507 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(112[14] 131[12])
    defparam period_counter__i7.GSR = "ENABLED";
    FD1S3IX period_counter__i6 (.D(period_counter_15__N_4409[6]), .CK(us_clk), 
            .CD(high_counter_9__N_4408), .Q(period_counter[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=19, LSE_RCOL=25, LSE_LLINE=495, LSE_RLINE=507 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(112[14] 131[12])
    defparam period_counter__i6.GSR = "ENABLED";
    FD1S3IX period_counter__i5 (.D(period_counter_15__N_4409[5]), .CK(us_clk), 
            .CD(high_counter_9__N_4408), .Q(period_counter[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=19, LSE_RCOL=25, LSE_LLINE=495, LSE_RLINE=507 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(112[14] 131[12])
    defparam period_counter__i5.GSR = "ENABLED";
    FD1S3IX period_counter__i4 (.D(n1[4]), .CK(us_clk), .CD(n30656), .Q(period_counter[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=19, LSE_RCOL=25, LSE_LLINE=495, LSE_RLINE=507 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(112[14] 131[12])
    defparam period_counter__i4.GSR = "ENABLED";
    FD1S3IX period_counter__i3 (.D(period_counter_15__N_4409[3]), .CK(us_clk), 
            .CD(high_counter_9__N_4408), .Q(period_counter[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=19, LSE_RCOL=25, LSE_LLINE=495, LSE_RLINE=507 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(112[14] 131[12])
    defparam period_counter__i3.GSR = "ENABLED";
    FD1S3IX period_counter__i2 (.D(n1[2]), .CK(us_clk), .CD(n30656), .Q(period_counter[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=19, LSE_RCOL=25, LSE_LLINE=495, LSE_RLINE=507 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(112[14] 131[12])
    defparam period_counter__i2.GSR = "ENABLED";
    FD1S3IX period_counter__i1 (.D(n1[1]), .CK(us_clk), .CD(n30656), .Q(period_counter[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=19, LSE_RCOL=25, LSE_LLINE=495, LSE_RLINE=507 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(112[14] 131[12])
    defparam period_counter__i1.GSR = "ENABLED";
    LUT4 i25766_2_lut (.A(n1[0]), .B(\next_state_2__N_4443[0] ), .Z(period_counter_15__N_4409[0])) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(127[14] 131[12])
    defparam i25766_2_lut.init = 16'heeee;
    CCU2D add_8_10 (.A0(high_counter[8]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(high_counter[9]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43819), .S0(n29[8]), .S1(n29[9]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(130[33:54])
    defparam add_8_10.INIT0 = 16'h5aaa;
    defparam add_8_10.INIT1 = 16'h5aaa;
    defparam add_8_10.INJECT1_0 = "NO";
    defparam add_8_10.INJECT1_1 = "NO";
    CCU2D add_8_8 (.A0(high_counter[6]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(high_counter[7]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n43818), .COUT(n43819), .S0(n29[6]), .S1(n29[7]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(130[33:54])
    defparam add_8_8.INIT0 = 16'h5aaa;
    defparam add_8_8.INIT1 = 16'h5aaa;
    defparam add_8_8.INJECT1_0 = "NO";
    defparam add_8_8.INJECT1_1 = "NO";
    FD1P3IX high_counter__i9 (.D(n29[9]), .SP(us_clk_enable_61), .CD(high_counter_9__N_4408), 
            .CK(us_clk), .Q(high_counter[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=19, LSE_RCOL=25, LSE_LLINE=495, LSE_RLINE=507 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(112[14] 131[12])
    defparam high_counter__i9.GSR = "ENABLED";
    CCU2D add_8_6 (.A0(high_counter[4]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(high_counter[5]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n43817), .COUT(n43818), .S0(n29[4]), .S1(n29[5]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(130[33:54])
    defparam add_8_6.INIT0 = 16'h5aaa;
    defparam add_8_6.INIT1 = 16'h5aaa;
    defparam add_8_6.INJECT1_0 = "NO";
    defparam add_8_6.INJECT1_1 = "NO";
    FD1P3IX high_counter__i8 (.D(n29[8]), .SP(us_clk_enable_61), .CD(high_counter_9__N_4408), 
            .CK(us_clk), .Q(high_counter[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=19, LSE_RCOL=25, LSE_LLINE=495, LSE_RLINE=507 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(112[14] 131[12])
    defparam high_counter__i8.GSR = "ENABLED";
    FD1P3IX high_counter__i7 (.D(n29[7]), .SP(us_clk_enable_61), .CD(high_counter_9__N_4408), 
            .CK(us_clk), .Q(high_counter[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=19, LSE_RCOL=25, LSE_LLINE=495, LSE_RLINE=507 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(112[14] 131[12])
    defparam high_counter__i7.GSR = "ENABLED";
    FD1P3IX high_counter__i6 (.D(n29[6]), .SP(us_clk_enable_61), .CD(high_counter_9__N_4408), 
            .CK(us_clk), .Q(high_counter[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=19, LSE_RCOL=25, LSE_LLINE=495, LSE_RLINE=507 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(112[14] 131[12])
    defparam high_counter__i6.GSR = "ENABLED";
    FD1P3IX high_counter__i5 (.D(n29[5]), .SP(us_clk_enable_61), .CD(high_counter_9__N_4408), 
            .CK(us_clk), .Q(high_counter[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=19, LSE_RCOL=25, LSE_LLINE=495, LSE_RLINE=507 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(112[14] 131[12])
    defparam high_counter__i5.GSR = "ENABLED";
    FD1P3IX high_counter__i4 (.D(n29[4]), .SP(us_clk_enable_61), .CD(high_counter_9__N_4408), 
            .CK(us_clk), .Q(high_counter[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=19, LSE_RCOL=25, LSE_LLINE=495, LSE_RLINE=507 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(112[14] 131[12])
    defparam high_counter__i4.GSR = "ENABLED";
    FD1P3IX high_counter__i3 (.D(n29[3]), .SP(us_clk_enable_61), .CD(high_counter_9__N_4408), 
            .CK(us_clk), .Q(high_counter[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=19, LSE_RCOL=25, LSE_LLINE=495, LSE_RLINE=507 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(112[14] 131[12])
    defparam high_counter__i3.GSR = "ENABLED";
    FD1P3IX high_counter__i2 (.D(n29[2]), .SP(us_clk_enable_61), .CD(high_counter_9__N_4408), 
            .CK(us_clk), .Q(high_counter[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=19, LSE_RCOL=25, LSE_LLINE=495, LSE_RLINE=507 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(112[14] 131[12])
    defparam high_counter__i2.GSR = "ENABLED";
    FD1P3IX high_counter__i1 (.D(n29[1]), .SP(us_clk_enable_61), .CD(high_counter_9__N_4408), 
            .CK(us_clk), .Q(high_counter[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=19, LSE_RCOL=25, LSE_LLINE=495, LSE_RLINE=507 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(112[14] 131[12])
    defparam high_counter__i1.GSR = "ENABLED";
    CCU2D add_8_4 (.A0(high_counter[2]), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(high_counter[3]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n43816), .COUT(n43817), .S0(n29[2]), .S1(n29[3]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(130[33:54])
    defparam add_8_4.INIT0 = 16'h5aaa;
    defparam add_8_4.INIT1 = 16'h5aaa;
    defparam add_8_4.INJECT1_0 = "NO";
    defparam add_8_4.INJECT1_1 = "NO";
    LUT4 i39658_2_lut (.A(\next_state_2__N_4443[0] ), .B(high_counter_9__N_4408), 
         .Z(n30656)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(112[14] 131[12])
    defparam i39658_2_lut.init = 16'heeee;
    CCU2D add_8_2 (.A0(high_counter[0]), .B0(high_counter_en), .C0(GND_net), 
          .D0(GND_net), .A1(high_counter[1]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n43816), .S1(n29[1]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(130[33:54])
    defparam add_8_2.INIT0 = 16'h7000;
    defparam add_8_2.INIT1 = 16'h5aaa;
    defparam add_8_2.INJECT1_0 = "NO";
    defparam add_8_2.INJECT1_1 = "NO";
    LUT4 i26269_2_lut (.A(n1[9]), .B(\next_state_2__N_4443[0] ), .Z(period_counter_15__N_4409[9])) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(127[14] 131[12])
    defparam i26269_2_lut.init = 16'heeee;
    LUT4 i26272_2_lut (.A(n1[8]), .B(\next_state_2__N_4443[0] ), .Z(period_counter_15__N_4409[8])) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(127[14] 131[12])
    defparam i26272_2_lut.init = 16'heeee;
    LUT4 i26275_2_lut (.A(n1[7]), .B(\next_state_2__N_4443[0] ), .Z(period_counter_15__N_4409[7])) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(127[14] 131[12])
    defparam i26275_2_lut.init = 16'heeee;
    LUT4 i26276_2_lut (.A(n1[6]), .B(\next_state_2__N_4443[0] ), .Z(period_counter_15__N_4409[6])) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(127[14] 131[12])
    defparam i26276_2_lut.init = 16'heeee;
    LUT4 i26277_2_lut (.A(n1[5]), .B(\next_state_2__N_4443[0] ), .Z(period_counter_15__N_4409[5])) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(127[14] 131[12])
    defparam i26277_2_lut.init = 16'heeee;
    LUT4 i26279_2_lut (.A(n1[3]), .B(\next_state_2__N_4443[0] ), .Z(period_counter_15__N_4409[3])) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(127[14] 131[12])
    defparam i26279_2_lut.init = 16'heeee;
    LUT4 i3_3_lut (.A(period_counter[4]), .B(period_counter[5]), .C(n27989), 
         .Z(n8)) /* synthesis lut_function=((B+(C))+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(112[18:50])
    defparam i3_3_lut.init = 16'hfdfd;
    LUT4 i39744_4_lut (.A(n27989), .B(n14_adj_5175), .C(n10), .D(period_counter[6]), 
         .Z(high_counter_9__N_4408)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(112[18:50])
    defparam i39744_4_lut.init = 16'h0001;
    LUT4 i6_4_lut (.A(period_counter[8]), .B(period_counter[7]), .C(n52406), 
         .D(period_counter[11]), .Z(n14_adj_5175)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;
    defparam i6_4_lut.init = 16'hfeff;
    LUT4 i33203_2_lut (.A(high_counter[0]), .B(high_counter_en), .Z(n29[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i33203_2_lut.init = 16'h6666;
    LUT4 i6_4_lut_adj_249 (.A(n11), .B(n9), .C(period_counter[0]), .D(period_counter[9]), 
         .Z(n27989)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(112[18:50])
    defparam i6_4_lut_adj_249.init = 16'hfeff;
    LUT4 i4_3_lut (.A(period_counter[2]), .B(period_counter[13]), .C(period_counter[12]), 
         .Z(n11)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(112[18:50])
    defparam i4_3_lut.init = 16'hfefe;
    LUT4 i2_2_lut (.A(period_counter[1]), .B(period_counter[15]), .Z(n9)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(112[18:50])
    defparam i2_2_lut.init = 16'heeee;
    CCU2D add_7_17 (.A0(period_counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n43814), .S0(n1[15]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(128[33:54])
    defparam add_7_17.INIT0 = 16'h5aaa;
    defparam add_7_17.INIT1 = 16'h0000;
    defparam add_7_17.INJECT1_0 = "NO";
    defparam add_7_17.INJECT1_1 = "NO";
    LUT4 i39689_4_lut (.A(n7), .B(period_counter[3]), .C(period_counter[10]), 
         .D(n27989), .Z(\next_state_2__N_4443[0] )) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(123[18:57])
    defparam i39689_4_lut.init = 16'h0004;
    LUT4 i4_4_lut (.A(n7_adj_5176), .B(period_counter[7]), .C(period_counter[8]), 
         .D(period_counter[14]), .Z(n47352)) /* synthesis lut_function=(A+(((D)+!C)+!B)) */ ;
    defparam i4_4_lut.init = 16'hffbf;
    LUT4 i2_2_lut_adj_250 (.A(period_counter[11]), .B(period_counter[6]), 
         .Z(n7_adj_5176)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i2_2_lut_adj_250.init = 16'hbbbb;
    LUT4 i1_2_lut_rep_469 (.A(period_counter[3]), .B(period_counter[10]), 
         .Z(n52405)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(112[18:50])
    defparam i1_2_lut_rep_469.init = 16'hbbbb;
    LUT4 i2_2_lut_3_lut (.A(period_counter[3]), .B(period_counter[10]), 
         .C(period_counter[14]), .Z(n10)) /* synthesis lut_function=(A+!(B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(112[18:50])
    defparam i2_2_lut_3_lut.init = 16'hbfbf;
    LUT4 i1_2_lut_rep_470 (.A(period_counter[4]), .B(period_counter[5]), 
         .Z(n52406)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(112[18:50])
    defparam i1_2_lut_rep_470.init = 16'hbbbb;
    LUT4 i2_2_lut_3_lut_adj_251 (.A(period_counter[4]), .B(period_counter[5]), 
         .C(n47352), .Z(n7)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(112[18:50])
    defparam i2_2_lut_3_lut_adj_251.init = 16'hfbfb;
    CCU2D add_7_15 (.A0(period_counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(period_counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43813), .COUT(n43814), .S0(n1[13]), .S1(n1[14]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(128[33:54])
    defparam add_7_15.INIT0 = 16'h5aaa;
    defparam add_7_15.INIT1 = 16'h5aaa;
    defparam add_7_15.INJECT1_0 = "NO";
    defparam add_7_15.INJECT1_1 = "NO";
    CCU2D add_7_13 (.A0(period_counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(period_counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43812), .COUT(n43813), .S0(n1[11]), .S1(n1[12]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(128[33:54])
    defparam add_7_13.INIT0 = 16'h5aaa;
    defparam add_7_13.INIT1 = 16'h5aaa;
    defparam add_7_13.INJECT1_0 = "NO";
    defparam add_7_13.INJECT1_1 = "NO";
    CCU2D add_7_11 (.A0(period_counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(period_counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43811), .COUT(n43812), .S0(n1[9]), .S1(n1[10]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(128[33:54])
    defparam add_7_11.INIT0 = 16'h5aaa;
    defparam add_7_11.INIT1 = 16'h5aaa;
    defparam add_7_11.INJECT1_0 = "NO";
    defparam add_7_11.INJECT1_1 = "NO";
    CCU2D add_7_9 (.A0(period_counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(period_counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43810), .COUT(n43811), .S0(n1[7]), .S1(n1[8]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(128[33:54])
    defparam add_7_9.INIT0 = 16'h5aaa;
    defparam add_7_9.INIT1 = 16'h5aaa;
    defparam add_7_9.INJECT1_0 = "NO";
    defparam add_7_9.INJECT1_1 = "NO";
    CCU2D add_7_7 (.A0(period_counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(period_counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43809), .COUT(n43810), .S0(n1[5]), .S1(n1[6]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(128[33:54])
    defparam add_7_7.INIT0 = 16'h5aaa;
    defparam add_7_7.INIT1 = 16'h5aaa;
    defparam add_7_7.INJECT1_0 = "NO";
    defparam add_7_7.INJECT1_1 = "NO";
    CCU2D add_7_5 (.A0(period_counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(period_counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43808), .COUT(n43809), .S0(n1[3]), .S1(n1[4]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(128[33:54])
    defparam add_7_5.INIT0 = 16'h5aaa;
    defparam add_7_5.INIT1 = 16'h5aaa;
    defparam add_7_5.INJECT1_0 = "NO";
    defparam add_7_5.INJECT1_1 = "NO";
    CCU2D add_7_3 (.A0(period_counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(period_counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43807), .COUT(n43808), .S0(n1[1]), .S1(n1[2]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(128[33:54])
    defparam add_7_3.INIT0 = 16'h5aaa;
    defparam add_7_3.INIT1 = 16'h5aaa;
    defparam add_7_3.INJECT1_0 = "NO";
    defparam add_7_3.INJECT1_1 = "NO";
    CCU2D add_7_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(period_counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n43807), .S1(n1[0]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(128[33:54])
    defparam add_7_1.INIT0 = 16'hF000;
    defparam add_7_1.INIT1 = 16'h5555;
    defparam add_7_1.INJECT1_0 = "NO";
    defparam add_7_1.INJECT1_1 = "NO";
    FD1P3IX high_counter_en_28 (.D(n53885), .SP(\next_state_2__N_4443[0] ), 
            .CD(high_counter_9__N_4408), .CK(us_clk), .Q(high_counter_en)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=19, LSE_RCOL=25, LSE_LLINE=495, LSE_RLINE=507 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(112[14] 131[12])
    defparam high_counter_en_28.GSR = "ENABLED";
    FD1S3IX period_counter__i15 (.D(n1[15]), .CK(us_clk), .CD(n30656), 
            .Q(period_counter[15])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=19, LSE_RCOL=25, LSE_LLINE=495, LSE_RLINE=507 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(112[14] 131[12])
    defparam period_counter__i15.GSR = "ENABLED";
    pwm_generator_block pwm4 (.\next_state_2__N_4440[2] (next_state_2__N_4440[2]), 
            .n48020(n48020), .resetn(resetn), .motor_4_pwm_c(motor_4_pwm_c), 
            .n36457(n36457), .\next_state_2__N_4443[0] (\next_state_2__N_4443[0] ), 
            .us_clk(us_clk), .high_counter_9__N_4408(high_counter_9__N_4408)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(89[25] 97[25])
    pwm_generator_block_U7 pwm3 (.n48749(n48749), .high_counter({high_counter}), 
            .\next_state_2__N_4440[2] (next_state_2__N_4440[2]), .n48020(n48020), 
            .resetn(resetn), .motor_3_pwm_c(motor_3_pwm_c), .n36457(n36457), 
            .\next_state_2__N_4443[0] (\next_state_2__N_4443[0] ), .us_clk(us_clk), 
            .high_counter_9__N_4408(high_counter_9__N_4408)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(78[25] 86[25])
    pwm_generator_block_U8 pwm2 (.resetn(resetn), .n36457(n36457), .n48020(n48020), 
            .\next_state_2__N_4440[2] (next_state_2__N_4440[2]), .motor_2_pwm_c(motor_2_pwm_c), 
            .\next_state_2__N_4443[0] (\next_state_2__N_4443[0] ), .us_clk(us_clk), 
            .high_counter_9__N_4408(high_counter_9__N_4408)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(67[25] 75[25])
    pwm_generator_block_U9 pwm1 (.\next_state_2__N_4440[2] (next_state_2__N_4440[2]), 
            .n48020(n48020), .resetn(resetn), .high_counter_9__N_4408(high_counter_9__N_4408), 
            .n48749(n48749), .n47352(n47352), .n8(n8), .n52405(n52405), 
            .n36457(n36457), .motor_1_pwm_c(motor_1_pwm_c), .\next_state_2__N_4443[0] (\next_state_2__N_4443[0] ), 
            .us_clk(us_clk)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator.v(56[25] 64[25])
    
endmodule
//
// Verilog Description of module pwm_generator_block
//

module pwm_generator_block (\next_state_2__N_4440[2] , n48020, resetn, 
            motor_4_pwm_c, n36457, \next_state_2__N_4443[0] , us_clk, 
            high_counter_9__N_4408) /* synthesis syn_module_defined=1 */ ;
    input \next_state_2__N_4440[2] ;
    input n48020;
    input resetn;
    output motor_4_pwm_c;
    input n36457;
    input \next_state_2__N_4443[0] ;
    input us_clk;
    input high_counter_9__N_4408;
    
    wire us_clk /* synthesis SET_AS_NETWORK=us_clk, is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(221[10:16])
    wire [2:0]state;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(44[15:20])
    wire [2:0]n10455;
    
    wire n10464, n48008, n26078, n36753, n5;
    
    LUT4 mux_4645_i3_4_lut (.A(state[0]), .B(\next_state_2__N_4440[2] ), 
         .C(state[2]), .D(n48020), .Z(n10455[2])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(56[9] 79[16])
    defparam mux_4645_i3_4_lut.init = 16'hc5c0;
    LUT4 i24_4_lut_3_lut (.A(state[1]), .B(state[0]), .C(state[2]), .Z(n10464)) /* synthesis lut_function=(A (B+(C))+!A (B (C)+!B !(C))) */ ;
    defparam i24_4_lut_3_lut.init = 16'he9e9;
    LUT4 i1_3_lut_4_lut (.A(resetn), .B(state[2]), .C(state[1]), .D(state[0]), 
         .Z(motor_4_pwm_c)) /* synthesis lut_function=(!((B+(C (D)+!C !(D)))+!A)) */ ;
    defparam i1_3_lut_4_lut.init = 16'h0220;
    LUT4 i39889_3_lut_4_lut (.A(resetn), .B(state[2]), .C(state[1]), .D(state[0]), 
         .Z(n48008)) /* synthesis lut_function=((B+(C (D)+!C !(D)))+!A) */ ;
    defparam i39889_3_lut_4_lut.init = 16'hfddf;
    LUT4 i14448_3_lut (.A(n36457), .B(\next_state_2__N_4443[0] ), .C(state[0]), 
         .Z(n26078)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(56[9] 79[16])
    defparam i14448_3_lut.init = 16'hcaca;
    FD1S3IX state_i2 (.D(n10455[2]), .CK(us_clk), .CD(n10464), .Q(state[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=25, LSE_RCOL=25, LSE_LLINE=89, LSE_RLINE=97 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(51[13:33])
    defparam state_i2.GSR = "ENABLED";
    LUT4 i39749_4_lut (.A(resetn), .B(n36753), .C(high_counter_9__N_4408), 
         .D(state[2]), .Z(n5)) /* synthesis lut_function=((B (C+!(D))+!B (C (D)))+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(56[9] 79[16])
    defparam i39749_4_lut.init = 16'hf5dd;
    LUT4 i26121_2_lut (.A(state[0]), .B(\next_state_2__N_4443[0] ), .Z(n36753)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(56[9] 79[16])
    defparam i26121_2_lut.init = 16'h2222;
    FD1S3IX state_i1 (.D(n26078), .CK(us_clk), .CD(n48008), .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=25, LSE_RCOL=25, LSE_LLINE=89, LSE_RLINE=97 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(51[13:33])
    defparam state_i1.GSR = "ENABLED";
    FD1S3JX state_i0 (.D(n5), .CK(us_clk), .PD(n10464), .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=25, LSE_RCOL=25, LSE_LLINE=89, LSE_RLINE=97 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(51[13:33])
    defparam state_i0.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module pwm_generator_block_U7
//

module pwm_generator_block_U7 (n48749, high_counter, \next_state_2__N_4440[2] , 
            n48020, resetn, motor_3_pwm_c, n36457, \next_state_2__N_4443[0] , 
            us_clk, high_counter_9__N_4408) /* synthesis syn_module_defined=1 */ ;
    output n48749;
    input [9:0]high_counter;
    input \next_state_2__N_4440[2] ;
    input n48020;
    input resetn;
    output motor_3_pwm_c;
    input n36457;
    input \next_state_2__N_4443[0] ;
    input us_clk;
    input high_counter_9__N_4408;
    
    wire us_clk /* synthesis SET_AS_NETWORK=us_clk, is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(221[10:16])
    
    wire n17, n15, n11, n12;
    wire [2:0]state;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(44[15:20])
    wire [2:0]n10428;
    
    wire n48005, n10437, n26073, n36761, n5;
    
    LUT4 i9_4_lut (.A(n17), .B(n15), .C(n11), .D(n12), .Z(n48749)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(68[26:53])
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 i7_4_lut (.A(high_counter[2]), .B(high_counter[8]), .C(high_counter[9]), 
         .D(high_counter[6]), .Z(n17)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(68[26:53])
    defparam i7_4_lut.init = 16'hfffe;
    LUT4 i5_2_lut (.A(high_counter[1]), .B(high_counter[5]), .Z(n15)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(68[26:53])
    defparam i5_2_lut.init = 16'heeee;
    LUT4 i1_2_lut (.A(high_counter[7]), .B(high_counter[4]), .Z(n11)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(68[26:53])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 i2_2_lut (.A(high_counter[0]), .B(high_counter[3]), .Z(n12)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(68[26:53])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 mux_4630_i3_4_lut (.A(state[0]), .B(\next_state_2__N_4440[2] ), 
         .C(state[2]), .D(n48020), .Z(n10428[2])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(56[9] 79[16])
    defparam mux_4630_i3_4_lut.init = 16'hc5c0;
    LUT4 i1_3_lut_4_lut (.A(resetn), .B(state[2]), .C(state[1]), .D(state[0]), 
         .Z(motor_3_pwm_c)) /* synthesis lut_function=(!((B+(C (D)+!C !(D)))+!A)) */ ;
    defparam i1_3_lut_4_lut.init = 16'h0220;
    LUT4 i39886_3_lut_4_lut (.A(resetn), .B(state[2]), .C(state[1]), .D(state[0]), 
         .Z(n48005)) /* synthesis lut_function=((B+(C (D)+!C !(D)))+!A) */ ;
    defparam i39886_3_lut_4_lut.init = 16'hfddf;
    LUT4 i24_4_lut_3_lut (.A(state[1]), .B(state[0]), .C(state[2]), .Z(n10437)) /* synthesis lut_function=(A (B+(C))+!A (B (C)+!B !(C))) */ ;
    defparam i24_4_lut_3_lut.init = 16'he9e9;
    LUT4 i14459_3_lut (.A(n36457), .B(\next_state_2__N_4443[0] ), .C(state[0]), 
         .Z(n26073)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(56[9] 79[16])
    defparam i14459_3_lut.init = 16'hcaca;
    FD1S3IX state_i2 (.D(n10428[2]), .CK(us_clk), .CD(n10437), .Q(state[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=25, LSE_RCOL=25, LSE_LLINE=78, LSE_RLINE=86 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(51[13:33])
    defparam state_i2.GSR = "ENABLED";
    LUT4 i39796_4_lut (.A(resetn), .B(n36761), .C(high_counter_9__N_4408), 
         .D(state[2]), .Z(n5)) /* synthesis lut_function=((B (C+!(D))+!B (C (D)))+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(56[9] 79[16])
    defparam i39796_4_lut.init = 16'hf5dd;
    LUT4 i26129_2_lut (.A(state[0]), .B(\next_state_2__N_4443[0] ), .Z(n36761)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(56[9] 79[16])
    defparam i26129_2_lut.init = 16'h2222;
    FD1S3IX state_i1 (.D(n26073), .CK(us_clk), .CD(n48005), .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=25, LSE_RCOL=25, LSE_LLINE=78, LSE_RLINE=86 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(51[13:33])
    defparam state_i1.GSR = "ENABLED";
    FD1S3JX state_i0 (.D(n5), .CK(us_clk), .PD(n10437), .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=25, LSE_RCOL=25, LSE_LLINE=78, LSE_RLINE=86 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(51[13:33])
    defparam state_i0.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module pwm_generator_block_U8
//

module pwm_generator_block_U8 (resetn, n36457, n48020, \next_state_2__N_4440[2] , 
            motor_2_pwm_c, \next_state_2__N_4443[0] , us_clk, high_counter_9__N_4408) /* synthesis syn_module_defined=1 */ ;
    input resetn;
    input n36457;
    output n48020;
    input \next_state_2__N_4440[2] ;
    output motor_2_pwm_c;
    input \next_state_2__N_4443[0] ;
    input us_clk;
    input high_counter_9__N_4408;
    
    wire us_clk /* synthesis SET_AS_NETWORK=us_clk, is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(221[10:16])
    wire [2:0]state;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(44[15:20])
    wire [2:0]n10401;
    
    wire n48002, n10410, n26068, n36767, n5;
    
    LUT4 i1_2_lut (.A(resetn), .B(n36457), .Z(n48020)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(56[9] 79[16])
    defparam i1_2_lut.init = 16'h2222;
    LUT4 mux_4615_i3_4_lut (.A(state[0]), .B(\next_state_2__N_4440[2] ), 
         .C(state[2]), .D(n48020), .Z(n10401[2])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(56[9] 79[16])
    defparam mux_4615_i3_4_lut.init = 16'hc5c0;
    LUT4 i1_3_lut_4_lut (.A(resetn), .B(state[2]), .C(state[1]), .D(state[0]), 
         .Z(motor_2_pwm_c)) /* synthesis lut_function=(!((B+(C (D)+!C !(D)))+!A)) */ ;
    defparam i1_3_lut_4_lut.init = 16'h0220;
    LUT4 i39883_3_lut_4_lut (.A(resetn), .B(state[2]), .C(state[1]), .D(state[0]), 
         .Z(n48002)) /* synthesis lut_function=((B+(C (D)+!C !(D)))+!A) */ ;
    defparam i39883_3_lut_4_lut.init = 16'hfddf;
    LUT4 i24_4_lut_3_lut (.A(state[1]), .B(state[0]), .C(state[2]), .Z(n10410)) /* synthesis lut_function=(A (B+(C))+!A (B (C)+!B !(C))) */ ;
    defparam i24_4_lut_3_lut.init = 16'he9e9;
    LUT4 i14480_3_lut (.A(n36457), .B(\next_state_2__N_4443[0] ), .C(state[0]), 
         .Z(n26068)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(56[9] 79[16])
    defparam i14480_3_lut.init = 16'hcaca;
    FD1S3IX state_i2 (.D(n10401[2]), .CK(us_clk), .CD(n10410), .Q(state[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=25, LSE_RCOL=25, LSE_LLINE=67, LSE_RLINE=75 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(51[13:33])
    defparam state_i2.GSR = "ENABLED";
    LUT4 i39787_4_lut (.A(resetn), .B(n36767), .C(high_counter_9__N_4408), 
         .D(state[2]), .Z(n5)) /* synthesis lut_function=((B (C+!(D))+!B (C (D)))+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(56[9] 79[16])
    defparam i39787_4_lut.init = 16'hf5dd;
    LUT4 i26135_2_lut (.A(state[0]), .B(\next_state_2__N_4443[0] ), .Z(n36767)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(56[9] 79[16])
    defparam i26135_2_lut.init = 16'h2222;
    FD1S3IX state_i1 (.D(n26068), .CK(us_clk), .CD(n48002), .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=25, LSE_RCOL=25, LSE_LLINE=67, LSE_RLINE=75 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(51[13:33])
    defparam state_i1.GSR = "ENABLED";
    FD1S3JX state_i0 (.D(n5), .CK(us_clk), .PD(n10410), .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=25, LSE_RCOL=25, LSE_LLINE=67, LSE_RLINE=75 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(51[13:33])
    defparam state_i0.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module pwm_generator_block_U9
//

module pwm_generator_block_U9 (\next_state_2__N_4440[2] , n48020, resetn, 
            high_counter_9__N_4408, n48749, n47352, n8, n52405, n36457, 
            motor_1_pwm_c, \next_state_2__N_4443[0] , us_clk) /* synthesis syn_module_defined=1 */ ;
    output \next_state_2__N_4440[2] ;
    input n48020;
    input resetn;
    input high_counter_9__N_4408;
    input n48749;
    input n47352;
    input n8;
    input n52405;
    output n36457;
    output motor_1_pwm_c;
    input \next_state_2__N_4443[0] ;
    input us_clk;
    
    wire us_clk /* synthesis SET_AS_NETWORK=us_clk, is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(221[10:16])
    wire [2:0]state;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(44[15:20])
    
    wire n10383;
    wire [2:0]n10374;
    
    wire n47999, n26063, n36773, n5;
    
    LUT4 i24_4_lut_3_lut (.A(state[1]), .B(state[0]), .C(state[2]), .Z(n10383)) /* synthesis lut_function=(A (B+(C))+!A (B (C)+!B !(C))) */ ;
    defparam i24_4_lut_3_lut.init = 16'he9e9;
    LUT4 mux_4600_i3_4_lut (.A(state[0]), .B(\next_state_2__N_4440[2] ), 
         .C(state[2]), .D(n48020), .Z(n10374[2])) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(56[9] 79[16])
    defparam mux_4600_i3_4_lut.init = 16'hc5c0;
    LUT4 i25837_2_lut (.A(resetn), .B(high_counter_9__N_4408), .Z(\next_state_2__N_4440[2] )) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam i25837_2_lut.init = 16'h2222;
    LUT4 i25835_4_lut (.A(n48749), .B(n47352), .C(n8), .D(n52405), .Z(n36457)) /* synthesis lut_function=(A (B+(C+(D)))) */ ;
    defparam i25835_4_lut.init = 16'haaa8;
    LUT4 i1_3_lut_4_lut (.A(resetn), .B(state[2]), .C(state[1]), .D(state[0]), 
         .Z(motor_1_pwm_c)) /* synthesis lut_function=(!((B+(C (D)+!C !(D)))+!A)) */ ;
    defparam i1_3_lut_4_lut.init = 16'h0220;
    LUT4 i39880_3_lut_4_lut (.A(resetn), .B(state[2]), .C(state[1]), .D(state[0]), 
         .Z(n47999)) /* synthesis lut_function=((B+(C (D)+!C !(D)))+!A) */ ;
    defparam i39880_3_lut_4_lut.init = 16'hfddf;
    LUT4 i14509_3_lut (.A(n36457), .B(\next_state_2__N_4443[0] ), .C(state[0]), 
         .Z(n26063)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(56[9] 79[16])
    defparam i14509_3_lut.init = 16'hcaca;
    FD1S3IX state_i2 (.D(n10374[2]), .CK(us_clk), .CD(n10383), .Q(state[2])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=25, LSE_RCOL=25, LSE_LLINE=56, LSE_RLINE=64 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(51[13:33])
    defparam state_i2.GSR = "ENABLED";
    LUT4 i39928_4_lut (.A(resetn), .B(n36773), .C(high_counter_9__N_4408), 
         .D(state[2]), .Z(n5)) /* synthesis lut_function=((B (C+!(D))+!B (C (D)))+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(56[9] 79[16])
    defparam i39928_4_lut.init = 16'hf5dd;
    LUT4 i26141_2_lut (.A(state[0]), .B(\next_state_2__N_4443[0] ), .Z(n36773)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(56[9] 79[16])
    defparam i26141_2_lut.init = 16'h2222;
    FD1S3IX state_i1 (.D(n26063), .CK(us_clk), .CD(n47999), .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=25, LSE_RCOL=25, LSE_LLINE=56, LSE_RLINE=64 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(51[13:33])
    defparam state_i1.GSR = "ENABLED";
    FD1S3JX state_i0 (.D(n5), .CK(us_clk), .PD(n10383), .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=10, LSE_LCOL=25, LSE_RCOL=25, LSE_LLINE=56, LSE_RLINE=64 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/pwm_generator_block.v(51[13:33])
    defparam state_i0.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module yaw_angle_accumulator
//

module yaw_angle_accumulator (n52179, \state[5] , \state[6] , n27995, 
            n37479) /* synthesis syn_module_defined=1 */ ;
    input n52179;
    input \state[5] ;
    input \state[6] ;
    input n27995;
    output n37479;
    
    
    LUT4 i26815_4_lut (.A(n52179), .B(\state[5] ), .C(\state[6] ), .D(n27995), 
         .Z(n37479)) /* synthesis lut_function=(A ((C+(D))+!B)) */ ;
    defparam i26815_4_lut.init = 16'haaa2;
    
endmodule
//
// Verilog Description of module \uart_top(NUM_DEBUG_ELEMENTS=8'b010010,FIXED_INTERVAL=0) 
//

module \uart_top(NUM_DEBUG_ELEMENTS=8'b010010,FIXED_INTERVAL=0)  (\tx_byte_index[0] , 
            \tx_byte_index[1] , n44797, swa_swb_val, n52359, \led_data[0] , 
            \led_data[3] , \led_data[2] , \led_data[1] , n50, n52, 
            VL53L1X_chip_id, n43303, n43217, \state[2] , n41683, \amc_debug[6] , 
            \amc_debug[5] , \state[5] , n52341, n52342, latched_pitch, 
            n15182, \z_linear_velocity[10] , \z_linear_velocity[8] , \z_linear_velocity[9] , 
            \z_linear_velocity[11] , sys_clk, \next_state[0] , \tx_word_index[1] , 
            VL53L1X_firm_rdy, throttle_val, n49177, \amc_debug[3] , 
            \amc_debug[2] , \amc_debug[1] , \amc_debug[7] , \VL53L1X_range_mm[9] , 
            \VL53L1X_range_mm[11] , \VL53L1X_range_mm[10] , \VL53L1X_range_mm[15] , 
            \VL53L1X_range_mm[14] , \VL53L1X_range_mm[13] , \z_linear_velocity[13] , 
            \z_linear_velocity[15] , \z_linear_velocity[14] , n48813, 
            n52441, n52456, yaw_val, n34690, n34692, \latched_roll[2] , 
            \state[6] , \VL53L1X_range_mm[4] , \VL53L1X_range_mm[7] , 
            \VL53L1X_range_mm[6] , \VL53L1X_range_mm[5] , n43332, n43302, 
            \z_linear_velocity[7] , \z_linear_velocity[4] , \z_linear_velocity[6] , 
            \z_linear_velocity[5] , \latched_roll[5] , \latched_roll[7] , 
            \latched_roll[6] , \VL53L1X_range_mm[12] , \z_linear_velocity[12] , 
            n44, n37479, \led_data[4] , n52179, n37731, n1406, n27995, 
            n38, \z_linear_velocity[3] , \z_linear_velocity[2] , \z_linear_velocity[1] , 
            n34474, VL53L1X_data_rdy, n43386, n34665, n51335, \latched_roll[4] , 
            \amc_debug[4] , \amc_debug[8] , n48820, GND_net, n52092, 
            n27, resetn_derived_2, n51271, n51272, n43221, n43225, 
            n10, \amc_debug[0] , n43309, n48081, n48828, n49185, 
            n52267, n52328, txrdy_n_c_7, n52255, n27734, \VL53L1X_range_mm[8] , 
            n51044, n52095, n51041, n123, n43271, n52390, n51201, 
            n51202, n51159, \i2c_device_driver_return_state[4] , n51273, 
            \VL53L1X_range_mm[1] , \VL53L1X_range_mm[2] , n52388, n52389, 
            n41688, n52429, n36752, n50674, n51135, n50715, n25, 
            n64, \led_data_out_7__N_1[2] , n50881, n52168, n52169, 
            \i2c_device_driver_return_state[0] , \i2c_device_driver_return_state[3] , 
            n52457, \next_dat_i_15__N_4452[3] , \next_state_4__N_1567[2] , 
            sout_c, sin_c, n53885, rxrdy_n_c, n53884) /* synthesis syn_module_defined=1 */ ;
    output \tx_byte_index[0] ;
    output \tx_byte_index[1] ;
    output n44797;
    input [7:0]swa_swb_val;
    output n52359;
    input \led_data[0] ;
    input \led_data[3] ;
    input \led_data[2] ;
    input \led_data[1] ;
    input n50;
    input n52;
    input [15:0]VL53L1X_chip_id;
    input n43303;
    input n43217;
    output \state[2] ;
    input n41683;
    input \amc_debug[6] ;
    input \amc_debug[5] ;
    output \state[5] ;
    output n52341;
    output n52342;
    input [7:0]latched_pitch;
    input n15182;
    input \z_linear_velocity[10] ;
    input \z_linear_velocity[8] ;
    input \z_linear_velocity[9] ;
    input \z_linear_velocity[11] ;
    input sys_clk;
    input \next_state[0] ;
    output \tx_word_index[1] ;
    input [7:0]VL53L1X_firm_rdy;
    input [7:0]throttle_val;
    input n49177;
    input \amc_debug[3] ;
    input \amc_debug[2] ;
    input \amc_debug[1] ;
    input \amc_debug[7] ;
    input \VL53L1X_range_mm[9] ;
    input \VL53L1X_range_mm[11] ;
    input \VL53L1X_range_mm[10] ;
    input \VL53L1X_range_mm[15] ;
    input \VL53L1X_range_mm[14] ;
    input \VL53L1X_range_mm[13] ;
    input \z_linear_velocity[13] ;
    input \z_linear_velocity[15] ;
    input \z_linear_velocity[14] ;
    input n48813;
    input n52441;
    input n52456;
    input [7:0]yaw_val;
    input n34690;
    input n34692;
    input \latched_roll[2] ;
    output \state[6] ;
    input \VL53L1X_range_mm[4] ;
    input \VL53L1X_range_mm[7] ;
    input \VL53L1X_range_mm[6] ;
    input \VL53L1X_range_mm[5] ;
    input n43332;
    input n43302;
    input \z_linear_velocity[7] ;
    input \z_linear_velocity[4] ;
    input \z_linear_velocity[6] ;
    input \z_linear_velocity[5] ;
    input \latched_roll[5] ;
    input \latched_roll[7] ;
    input \latched_roll[6] ;
    input \VL53L1X_range_mm[12] ;
    input \z_linear_velocity[12] ;
    output n44;
    input n37479;
    input \led_data[4] ;
    output n52179;
    output n37731;
    input n1406;
    output n27995;
    input n38;
    input \z_linear_velocity[3] ;
    input \z_linear_velocity[2] ;
    input \z_linear_velocity[1] ;
    input n34474;
    input [7:0]VL53L1X_data_rdy;
    input n43386;
    input n34665;
    input n51335;
    input \latched_roll[4] ;
    input \amc_debug[4] ;
    input \amc_debug[8] ;
    input n48820;
    input GND_net;
    input n52092;
    input n27;
    input resetn_derived_2;
    output n51271;
    output n51272;
    input n43221;
    input n43225;
    output n10;
    input \amc_debug[0] ;
    input n43309;
    output n48081;
    input n48828;
    input n49185;
    input n52267;
    output n52328;
    output txrdy_n_c_7;
    output n52255;
    output n27734;
    input \VL53L1X_range_mm[8] ;
    input n51044;
    input n52095;
    input n51041;
    output n123;
    input n43271;
    input n52390;
    input n51201;
    input n51202;
    input n51159;
    input \i2c_device_driver_return_state[4] ;
    input n51273;
    input \VL53L1X_range_mm[1] ;
    input \VL53L1X_range_mm[2] ;
    input n52388;
    input n52389;
    input n41688;
    input n52429;
    input n36752;
    input n50674;
    input n51135;
    input n50715;
    input n25;
    output n64;
    output \led_data_out_7__N_1[2] ;
    input n50881;
    input n52168;
    input n52169;
    input \i2c_device_driver_return_state[0] ;
    input \i2c_device_driver_return_state[3] ;
    input n52457;
    input \next_dat_i_15__N_4452[3] ;
    input \next_state_4__N_1567[2] ;
    output sout_c;
    input sin_c;
    input n53885;
    output rxrdy_n_c;
    input n53884;
    
    wire sys_clk /* synthesis SET_AS_NETWORK=sys_clk, is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(220[10:17])
    
    wire n3, n52530;
    wire [3:0]tx_byte_index;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(96[17:30])
    wire [15:0]n9499;
    
    wire n39, n34503, n34504, n18, n30, n1, n52158, n49377, 
        n51317, n51318, n48129, n52244, n7;
    wire [9:0]state;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(92[29:34])
    
    wire n25954, n25955, n48199, n49734, n49735;
    wire [7:0]tx_word_index;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(97[17:30])
    
    wire n49738, n49740, n1_adj_5106, n53077, n49736, n49737, n49739, 
        n50864, n51157, n27_c, n2, n47335, n52379, n50956, n4, 
        n52497, n52272, n47964, n47968, n52529, n52528, n38329, 
        n49424, n52532, n52453, n52451, n52258, n22;
    wire [9:0]next_state_9__N_4478;
    
    wire n38325, n49423, n52531, n52245, n52294, n44893, n52510, 
        n52511, n52512, n51327, next_state_9__N_4614, n49291, n13, 
        n27_adj_5107, n14, n27_adj_5108, n52184, n47346, n52178, 
        sys_clk_enable_246, n52541;
    wire [7:0]adr_i;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(87[29:34])
    wire [7:0]next_adr_i_7__N_4470;
    
    wire we_i, n52196, n51581, n51580, n34729, n52596, n3_adj_5109, 
        n52454, n51612, n52437, n51610, n51613, n51045, n2_adj_5110, 
        n3_adj_5111, n3_adj_5112, n11, n49484, n52562, n52561, n48861, 
        n51629, n52568, n52567, n50884, n1_adj_5113, n6, n48161, 
        n52141, n52586, n52585, n49448, n3_adj_5114, n53075, n52595, 
        n52594, n52598, n52597, n48147, n52143, n65, n89, n49, 
        n38081, n50897, n52398;
    wire [15:0]n9354;
    
    wire n24, n99, n38059, n50895, n50907, n27_adj_5115, n51009, 
        n51008, n53874, n23, n34534, n53235, n49411, n50860, n53233, 
        n53869, n52716, n53238, n53239, n53237, n53240, n51017, 
        n3_adj_5116, cyc_i;
    wire [9:0]next_state_9__N_4541;
    
    wire n38167, n53383, n49709, n51029, n49708, n51742, n48537, 
        n71, n6_adj_5117, n2_adj_5118, n49706, n51743, n53381, n14_adj_5119, 
        n51746, n51747, n38035, n53396, n53394, n50675, n20, n27_adj_5120, 
        n25_c, n40, n38267, n38447, n52206, n49281, n4_adj_5121, 
        n31, n48229, n49106, n22616, n53527;
    wire [15:0]n2019;
    
    wire n53525, n53523, n53524, n53559, n53558, n53557, n52208, 
        n50676, n51, n48706, n27_adj_5122, n22_adj_5123, n38023, 
        n50975, n50977, n52718, n51353, n52413, n26246, n27740, 
        n52587, n47966, n53870, n53776, n41729, n23_adj_5124, n52180, 
        n21, n49429, n52173, n49483, n49485, n52375, n38373, n52295, 
        n48742, n34493, n52207, n53773, n50859, n52443, n25919, 
        n91, n99_adj_5125, n47965, n13_adj_5126, n51016, n47969, 
        n51328, n47967, n52715, n13_adj_5127, n52166, n49376, n51326, 
        n13_adj_5128, n51336, n52164, n37957;
    wire [15:0]n1524;
    
    wire n21_adj_5129, n52434;
    wire [15:0]n304;
    
    wire n51324, n51323, n51325, n51027, n50807, n49381, n53398, 
        n51972, n51028, n53385, n51974, n50_adj_5130, n5, n7_adj_5131, 
        n51321, n50855, n51322, n51319, n51320, n48143, n38079, 
        n49482, n25965, n53076, n37942, n37950, n52165, n38458, 
        n121, n52717, n52496, n52495, n48679, n51316, n49426, 
        n49427, n52414, n47986, n52391, n52096, n43869;
    wire [7:0]n8;
    
    wire n49435, n43868, n50806, n50805, n52155, n48692, n19, 
        n37943, n37951, n37975, n52383;
    wire [3:0]n9;
    
    wire n43867;
    wire [15:0]dat_i;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(86[29:34])
    wire [15:0]next_dat_i_15__N_4452;
    
    wire n49682, n49431, n52395, n43866, n42210, n42214, n48839, 
        n52399, n52167, n52378, n50747, n50746, n52160, n49697, 
        n52407, n27651, n51047, n23_adj_5139, n50718, n50719, n5_adj_5140, 
        n6_adj_5141, n53078, n49085, n27742, n27743, n25959, n27741, 
        n51631, n48972, n48486, n48928, n48969, n49401, n47988, 
        n51975, n47990, n49712, n47989, n4_adj_5142, n52563, n52419, 
        n50720, n50721;
    wire [9:0]next_state_9__N_4551;
    
    wire n47985, n52599, sys_clk_enable_236, n38171, n14_adj_5144, 
        n52257, n14_adj_5145, n14_adj_5146, n47987, n52422, n51042, 
        n40166, n123_c, n86, n48589, n81, n85, n37, n49126, 
        n39_adj_5147;
    wire [9:0]next_state_9__N_4571;
    wire [9:0]next_state_9__N_4531;
    
    wire n20_adj_5148, n51046, n51043, n52097, n26269, n108, n117, 
        n41_adj_5149, n108_adj_5150, n117_adj_5151, n108_adj_5152, n117_adj_5153, 
        n108_adj_5155, n117_adj_5156, n123_adj_5157, n108_adj_5158, 
        n117_adj_5159;
    wire [15:0]n2147;
    
    wire n37965, n51289, n15, n3_adj_5160, n108_adj_5161, n117_adj_5162, 
        n17, n51351, n121_adj_5163, n51015, n53871, n25957, n48295, 
        n38452, n38456, n27735, n48731, n52240, n7_adj_5164, n47552, 
        n52442, n48676, n27_adj_5165, n12, n36607, n14_adj_5166, 
        n12_adj_5167, n50824, n22_adj_5168, n25927, n114, n6_adj_5169, 
        n38444, n38454, n45947, n4_adj_5170, n25964, n49476, n50858, 
        n48823, n28, n12_adj_5171, n51611, n51627, n51748, n51744, 
        n49710, n49711, n38432, n14_adj_5172, n50886, n49399, n49400, 
        n53526, n53397, n53395, n51749, n53384, n53382, n51745, 
        n52194, n52195, sys_clk_enable_217, n53236, n53234, n40212, 
        n50896, n6_adj_5174, n50882, n51630, n51628;
    
    LUT4 i39234_3_lut (.A(n3), .B(n52530), .C(tx_byte_index[2]), .Z(n9499[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(333[21] 354[28])
    defparam i39234_3_lut.init = 16'hcaca;
    PFUMX i23861 (.BLUT(n39), .ALUT(n34503), .C0(\tx_byte_index[0] ), 
          .Z(n34504));
    LUT4 i1_4_lut_4_lut_4_lut (.A(\tx_byte_index[1] ), .B(tx_byte_index[3]), 
         .C(tx_byte_index[2]), .D(n18), .Z(n30)) /* synthesis lut_function=(A (B+(C))+!A (B+!(C+!(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam i1_4_lut_4_lut_4_lut.init = 16'hedec;
    LUT4 i38582_3_lut_3_lut_4_lut (.A(tx_byte_index[2]), .B(\tx_byte_index[1] ), 
         .C(n1), .D(n52158), .Z(n49377)) /* synthesis lut_function=(A (D)+!A !(B+!(C))) */ ;
    defparam i38582_3_lut_3_lut_4_lut.init = 16'hba10;
    LUT4 n51317_bdd_3_lut_3_lut_4_lut (.A(tx_byte_index[2]), .B(\tx_byte_index[1] ), 
         .C(n1), .D(n51317), .Z(n51318)) /* synthesis lut_function=(A (D)+!A !(B+!(C))) */ ;
    defparam n51317_bdd_3_lut_3_lut_4_lut.init = 16'hba10;
    LUT4 i1_2_lut_3_lut_4_lut (.A(n48129), .B(n52244), .C(n7), .D(state[7]), 
         .Z(n44797)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B (C+!(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(366[17:29])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0f0e;
    LUT4 i1_2_lut_rep_423 (.A(swa_swb_val[2]), .B(swa_swb_val[1]), .Z(n52359)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i1_2_lut_rep_423.init = 16'heeee;
    LUT4 i15481_3_lut_4_lut (.A(\tx_byte_index[1] ), .B(n1), .C(n25954), 
         .D(tx_byte_index[2]), .Z(n25955)) /* synthesis lut_function=(A (C (D))+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(333[21] 354[28])
    defparam i15481_3_lut_4_lut.init = 16'hf044;
    LUT4 i1_2_lut_3_lut (.A(swa_swb_val[2]), .B(swa_swb_val[1]), .C(swa_swb_val[3]), 
         .Z(n48199)) /* synthesis lut_function=(A+(B+!(C))) */ ;
    defparam i1_2_lut_3_lut.init = 16'hefef;
    L6MUX21 i38943 (.D0(n49734), .D1(n49735), .SD(tx_word_index[0]), .Z(n49738));
    LUT4 n49448_bdd_4_lut (.A(n49740), .B(n1_adj_5106), .C(\tx_byte_index[1] ), 
         .D(tx_byte_index[2]), .Z(n53077)) /* synthesis lut_function=(A (B ((D)+!C)+!B (D))+!A !((C+(D))+!B)) */ ;
    defparam n49448_bdd_4_lut.init = 16'haa0c;
    L6MUX21 i38944 (.D0(n49736), .D1(n49737), .SD(tx_word_index[0]), .Z(n49739));
    LUT4 led_data_0__bdd_4_lut_41583 (.A(\led_data[0] ), .B(\led_data[3] ), 
         .C(\led_data[2] ), .D(\led_data[1] ), .Z(n50864)) /* synthesis lut_function=(!(A (B (C+(D)))+!A !(B (C+(D))))) */ ;
    defparam led_data_0__bdd_4_lut_41583.init = 16'h666a;
    LUT4 i1_4_lut (.A(\tx_byte_index[1] ), .B(swa_swb_val[0]), .C(n51157), 
         .D(swa_swb_val[3]), .Z(n27_c)) /* synthesis lut_function=(A+(B (C+!(D))+!B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(265[13] 275[20])
    defparam i1_4_lut.init = 16'hfaee;
    PFUMX i24154 (.BLUT(n50), .ALUT(n52), .C0(\tx_byte_index[0] ), .Z(n2));
    LUT4 n50955_bdd_2_lut_3_lut_4_lut (.A(tx_word_index[4]), .B(n47335), 
         .C(tx_word_index[2]), .D(n52379), .Z(n50956)) /* synthesis lut_function=(A+(B+(C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(335[25:29])
    defparam n50955_bdd_2_lut_3_lut_4_lut.init = 16'hfeee;
    LUT4 i1_2_lut_4_lut (.A(n4), .B(n52497), .C(n52272), .D(n47964), 
         .Z(n47968)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_2_lut_4_lut.init = 16'hca00;
    LUT4 n51845_bdd_4_lut_then_4_lut (.A(VL53L1X_chip_id[3]), .B(VL53L1X_chip_id[1]), 
         .C(\tx_byte_index[1] ), .D(VL53L1X_chip_id[2]), .Z(n52529)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (C)) */ ;
    defparam n51845_bdd_4_lut_then_4_lut.init = 16'hf0f2;
    LUT4 n51845_bdd_4_lut_else_4_lut (.A(VL53L1X_chip_id[5]), .B(\tx_byte_index[1] ), 
         .C(VL53L1X_chip_id[7]), .D(VL53L1X_chip_id[6]), .Z(n52528)) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;
    defparam n51845_bdd_4_lut_else_4_lut.init = 16'hccdc;
    LUT4 i38629_4_lut (.A(n38329), .B(\tx_byte_index[1] ), .C(tx_byte_index[2]), 
         .D(n43303), .Z(n49424)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;
    defparam i38629_4_lut.init = 16'hfaca;
    LUT4 i1_4_lut_4_lut_then_4_lut (.A(tx_byte_index[3]), .B(tx_word_index[2]), 
         .C(n47335), .D(tx_word_index[4]), .Z(n52532)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam i1_4_lut_4_lut_then_4_lut.init = 16'h0001;
    LUT4 i2_3_lut_4_lut (.A(n52453), .B(n52451), .C(n52258), .D(n22), 
         .Z(next_state_9__N_4478[1])) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i2_3_lut_4_lut.init = 16'h0100;
    LUT4 i38628_4_lut (.A(n38325), .B(\tx_byte_index[1] ), .C(tx_byte_index[2]), 
         .D(n43217), .Z(n49423)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;
    defparam i38628_4_lut.init = 16'hfaca;
    LUT4 i1_4_lut_4_lut_else_4_lut (.A(tx_byte_index[3]), .B(n47335), .C(tx_word_index[4]), 
         .Z(n52531)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam i1_4_lut_4_lut_else_4_lut.init = 16'h0101;
    LUT4 i1_3_lut_4_lut (.A(n52245), .B(n52294), .C(state[0]), .D(state[1]), 
         .Z(n44893)) /* synthesis lut_function=(!(A+(B+(C (D)+!C !(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(299[17:22])
    defparam i1_3_lut_4_lut.init = 16'h0110;
    PFUMX i40934 (.BLUT(n52510), .ALUT(n52511), .C0(\state[2] ), .Z(n52512));
    LUT4 n41683_bdd_4_lut (.A(n41683), .B(\amc_debug[6] ), .C(\amc_debug[5] ), 
         .D(\tx_byte_index[1] ), .Z(n51327)) /* synthesis lut_function=(A (C+(D))+!A (B ((D)+!C)+!B (D))) */ ;
    defparam n41683_bdd_4_lut.init = 16'hffa4;
    LUT4 i2_3_lut_4_lut_adj_149 (.A(n52245), .B(n52294), .C(state[0]), 
         .D(state[1]), .Z(next_state_9__N_4614)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(299[17:22])
    defparam i2_3_lut_4_lut_adj_149.init = 16'hffef;
    LUT4 i38499_2_lut_3_lut_4_lut (.A(\state[5] ), .B(n52341), .C(state[9]), 
         .D(n52342), .Z(n49291)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i38499_2_lut_3_lut_4_lut.init = 16'hfffe;
    PFUMX i38942 (.BLUT(n13), .ALUT(n27_adj_5107), .C0(\tx_byte_index[0] ), 
          .Z(n49737));
    LUT4 i1_4_lut_adj_150 (.A(\tx_byte_index[1] ), .B(latched_pitch[0]), 
         .C(n14), .D(latched_pitch[3]), .Z(n27_adj_5108)) /* synthesis lut_function=(A+(B (C+!(D))+!B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(265[13] 275[20])
    defparam i1_4_lut_adj_150.init = 16'hfaee;
    LUT4 i1_2_lut_4_lut_adj_151 (.A(n52184), .B(n47346), .C(n52178), .D(n15182), 
         .Z(sys_clk_enable_246)) /* synthesis lut_function=(A (B (D)+!B (C+(D)))+!A (D)) */ ;
    defparam i1_2_lut_4_lut_adj_151.init = 16'hff20;
    LUT4 tx_word_index_0__bdd_3_lut_then_4_lut (.A(\z_linear_velocity[10] ), 
         .B(\z_linear_velocity[8] ), .C(\z_linear_velocity[9] ), .D(\z_linear_velocity[11] ), 
         .Z(n52541)) /* synthesis lut_function=(A (B+(C+!(D)))) */ ;
    defparam tx_word_index_0__bdd_3_lut_then_4_lut.init = 16'ha8aa;
    FD1S3AX adr_i_i1 (.D(next_adr_i_7__N_4470[0]), .CK(sys_clk), .Q(adr_i[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=64, LSE_RCOL=6, LSE_LLINE=528, LSE_RLINE=562 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam adr_i_i1.GSR = "ENABLED";
    FD1S3AX state_i0 (.D(\next_state[0] ), .CK(sys_clk), .Q(state[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=64, LSE_RCOL=6, LSE_LLINE=528, LSE_RLINE=562 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam state_i0.GSR = "ENABLED";
    FD1S3AX we_i_417 (.D(next_state_9__N_4614), .CK(sys_clk), .Q(we_i)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=64, LSE_RCOL=6, LSE_LLINE=528, LSE_RLINE=562 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam we_i_417.GSR = "ENABLED";
    LUT4 i2_3_lut_rep_260_4_lut (.A(n52245), .B(n52294), .C(state[0]), 
         .D(state[1]), .Z(n52196)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(299[17:22])
    defparam i2_3_lut_rep_260_4_lut.init = 16'hfeff;
    LUT4 tx_word_index_3__bdd_4_lut (.A(tx_word_index[5]), .B(tx_word_index[4]), 
         .C(tx_word_index[7]), .D(tx_word_index[6]), .Z(n51581)) /* synthesis lut_function=(A (B+!(C))+!A !(B+!(C (D)))) */ ;
    defparam tx_word_index_3__bdd_4_lut.init = 16'h9a8a;
    LUT4 tx_word_index_3__bdd_4_lut_40529 (.A(tx_word_index[3]), .B(tx_word_index[2]), 
         .C(\tx_word_index[1] ), .D(tx_word_index[0]), .Z(n51580)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (C (D)))+!A (C)) */ ;
    defparam tx_word_index_3__bdd_4_lut_40529.init = 16'hf058;
    LUT4 i1_3_lut (.A(n34729), .B(\tx_byte_index[1] ), .C(n52596), .Z(n3_adj_5109)) /* synthesis lut_function=(A+(B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(96[17:30])
    defparam i1_3_lut.init = 16'heaea;
    LUT4 i2_3_lut_rep_248_4_lut (.A(n52454), .B(n52245), .C(state[4]), 
         .D(n52451), .Z(n52184)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam i2_3_lut_rep_248_4_lut.init = 16'hffef;
    LUT4 VL53L1X_firm_rdy_5__bdd_4_lut_40842 (.A(VL53L1X_firm_rdy[5]), .B(VL53L1X_firm_rdy[7]), 
         .C(VL53L1X_firm_rdy[4]), .D(VL53L1X_firm_rdy[6]), .Z(n51612)) /* synthesis lut_function=(A ((C)+!B)+!A !((C+!(D))+!B)) */ ;
    defparam VL53L1X_firm_rdy_5__bdd_4_lut_40842.init = 16'ha6a2;
    LUT4 i1_2_lut_rep_501 (.A(throttle_val[5]), .B(throttle_val[7]), .Z(n52437)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_rep_501.init = 16'hbbbb;
    LUT4 n11_bdd_4_lut_40638 (.A(VL53L1X_firm_rdy[1]), .B(VL53L1X_firm_rdy[3]), 
         .C(VL53L1X_firm_rdy[0]), .D(VL53L1X_firm_rdy[2]), .Z(n51610)) /* synthesis lut_function=(A ((C)+!B)+!A !((C+!(D))+!B)) */ ;
    defparam n11_bdd_4_lut_40638.init = 16'ha6a2;
    LUT4 n51612_bdd_2_lut (.A(n51612), .B(\tx_byte_index[1] ), .Z(n51613)) /* synthesis lut_function=(A+(B)) */ ;
    defparam n51612_bdd_2_lut.init = 16'heeee;
    LUT4 n48138_bdd_2_lut_40337_3_lut (.A(throttle_val[5]), .B(throttle_val[7]), 
         .C(throttle_val[6]), .Z(n51045)) /* synthesis lut_function=(A+((C)+!B)) */ ;
    defparam n48138_bdd_2_lut_40337_3_lut.init = 16'hfbfb;
    LUT4 i1_3_lut_adj_152 (.A(\tx_byte_index[1] ), .B(n34729), .C(n2_adj_5110), 
         .Z(n3_adj_5111)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(96[17:30])
    defparam i1_3_lut_adj_152.init = 16'hecec;
    PFUMX i38689 (.BLUT(n3_adj_5112), .ALUT(n11), .C0(\tx_byte_index[0] ), 
          .Z(n49484));
    LUT4 n60_bdd_4_lut_then_3_lut (.A(VL53L1X_chip_id[10]), .B(VL53L1X_chip_id[11]), 
         .C(VL53L1X_chip_id[9]), .Z(n52562)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam n60_bdd_4_lut_then_3_lut.init = 16'hc8c8;
    LUT4 n60_bdd_4_lut_else_3_lut (.A(VL53L1X_chip_id[13]), .B(VL53L1X_chip_id[15]), 
         .C(VL53L1X_chip_id[14]), .Z(n52561)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam n60_bdd_4_lut_else_3_lut.init = 16'hc8c8;
    LUT4 n9512_bdd_4_lut (.A(n34729), .B(\tx_byte_index[1] ), .C(tx_byte_index[2]), 
         .D(n48861), .Z(n51629)) /* synthesis lut_function=(A (B+!(C (D)))+!A (B (C)+!B !((D)+!C))) */ ;
    defparam n9512_bdd_4_lut.init = 16'hcafa;
    LUT4 i5_4_lut (.A(state[8]), .B(n52342), .C(n52341), .D(n52512), 
         .Z(next_state_9__N_4478[3])) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i5_4_lut.init = 16'h0100;
    LUT4 n300_bdd_4_lut_then_4_lut (.A(tx_word_index[3]), .B(\tx_word_index[1] ), 
         .C(\tx_byte_index[1] ), .D(tx_word_index[2]), .Z(n52568)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam n300_bdd_4_lut_then_4_lut.init = 16'h0002;
    LUT4 n300_bdd_4_lut_else_4_lut (.A(tx_word_index[5]), .B(\tx_byte_index[1] ), 
         .C(tx_word_index[6]), .D(tx_word_index[7]), .Z(n52567)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam n300_bdd_4_lut_else_4_lut.init = 16'h0100;
    LUT4 n48198_bdd_3_lut_40832 (.A(swa_swb_val[5]), .B(swa_swb_val[7]), 
         .C(swa_swb_val[6]), .Z(n50884)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam n48198_bdd_3_lut_40832.init = 16'hc8c8;
    PFUMX i25573 (.BLUT(n1_adj_5113), .ALUT(n6), .C0(\tx_byte_index[0] ), 
          .Z(n2_adj_5110));
    LUT4 VL53L1X_firm_rdy_2__bdd_4_lut_41589 (.A(VL53L1X_firm_rdy[2]), .B(n48161), 
         .C(n49177), .D(tx_word_index[0]), .Z(n52141)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam VL53L1X_firm_rdy_2__bdd_4_lut_41589.init = 16'hf011;
    LUT4 n48960_bdd_4_lut_then_4_lut (.A(\amc_debug[3] ), .B(\amc_debug[2] ), 
         .C(\tx_byte_index[1] ), .D(\amc_debug[1] ), .Z(n52586)) /* synthesis lut_function=(A (B (C)+!B (C+!(D)))+!A (C)) */ ;
    defparam n48960_bdd_4_lut_then_4_lut.init = 16'hf0f2;
    LUT4 n48960_bdd_4_lut_else_4_lut (.A(\amc_debug[5] ), .B(\tx_byte_index[1] ), 
         .C(\amc_debug[6] ), .D(\amc_debug[7] ), .Z(n52585)) /* synthesis lut_function=(A (B)+!A (B+!(C+!(D)))) */ ;
    defparam n48960_bdd_4_lut_else_4_lut.init = 16'hcdcc;
    LUT4 n49448_bdd_4_lut_41232 (.A(n49448), .B(n3_adj_5114), .C(tx_byte_index[2]), 
         .D(tx_word_index[0]), .Z(n53075)) /* synthesis lut_function=(A (B+(C+!(D)))+!A !((C+!(D))+!B)) */ ;
    defparam n49448_bdd_4_lut_41232.init = 16'hacaa;
    LUT4 VL53L1X_range_mm_15__bdd_4_lut_then_3_lut (.A(\VL53L1X_range_mm[9] ), 
         .B(\VL53L1X_range_mm[11] ), .C(\VL53L1X_range_mm[10] ), .Z(n52595)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam VL53L1X_range_mm_15__bdd_4_lut_then_3_lut.init = 16'h0404;
    LUT4 VL53L1X_range_mm_15__bdd_4_lut_else_3_lut (.A(\VL53L1X_range_mm[15] ), 
         .B(\VL53L1X_range_mm[14] ), .C(\VL53L1X_range_mm[13] ), .Z(n52594)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;
    defparam VL53L1X_range_mm_15__bdd_4_lut_else_3_lut.init = 16'h0202;
    LUT4 n14_bdd_4_lut_then_3_lut (.A(\z_linear_velocity[9] ), .B(\z_linear_velocity[11] ), 
         .C(\z_linear_velocity[10] ), .Z(n52598)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam n14_bdd_4_lut_then_3_lut.init = 16'hc8c8;
    LUT4 n14_bdd_4_lut_else_3_lut (.A(\z_linear_velocity[13] ), .B(\z_linear_velocity[15] ), 
         .C(\z_linear_velocity[14] ), .Z(n52597)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam n14_bdd_4_lut_else_3_lut.init = 16'hc8c8;
    LUT4 VL53L1X_firm_rdy_6__bdd_4_lut (.A(VL53L1X_firm_rdy[6]), .B(n48147), 
         .C(n48813), .D(tx_word_index[0]), .Z(n52143)) /* synthesis lut_function=(A (C (D))+!A (B (C (D))+!B (C+!(D)))) */ ;
    defparam VL53L1X_firm_rdy_6__bdd_4_lut.init = 16'hf011;
    PFUMX i42 (.BLUT(n65), .ALUT(n89), .C0(\tx_byte_index[0] ), .Z(n49));
    LUT4 n18_bdd_4_lut_40825 (.A(n38081), .B(n52441), .C(throttle_val[3]), 
         .D(\tx_byte_index[0] ), .Z(n50897)) /* synthesis lut_function=(A (B (C+!(D))+!B !(D))+!A (B (C (D)))) */ ;
    defparam n18_bdd_4_lut_40825.init = 16'hc0aa;
    LUT4 i39312_3_lut_4_lut_4_lut (.A(n52398), .B(n9354[6]), .C(tx_word_index[0]), 
         .D(n24), .Z(n99)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i39312_3_lut_4_lut_4_lut.init = 16'hc5c0;
    LUT4 n18_bdd_4_lut_40106 (.A(n38059), .B(n52456), .C(\tx_byte_index[0] ), 
         .D(yaw_val[3]), .Z(n50895)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;
    defparam n18_bdd_4_lut_40106.init = 16'hca0a;
    LUT4 n314_bdd_4_lut_40905 (.A(tx_word_index[4]), .B(tx_word_index[7]), 
         .C(tx_word_index[6]), .D(tx_word_index[5]), .Z(n50907)) /* synthesis lut_function=(!(A (B (C+(D)))+!A !(B (C+(D))))) */ ;
    defparam n314_bdd_4_lut_40905.init = 16'h666a;
    LUT4 i1_4_lut_adj_153 (.A(\tx_byte_index[1] ), .B(n34690), .C(n34692), 
         .D(\latched_roll[2] ), .Z(n27_adj_5115)) /* synthesis lut_function=(A+(B (C+!(D))+!B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(265[13] 275[20])
    defparam i1_4_lut_adj_153.init = 16'hfaee;
    LUT4 n51009_bdd_4_lut (.A(n51009), .B(n51008), .C(\tx_byte_index[0] ), 
         .D(\tx_byte_index[1] ), .Z(n53874)) /* synthesis lut_function=(!(A (B (C (D))+!B (C))+!A (B (C (D)+!C !(D))+!B (C+!(D))))) */ ;
    defparam n51009_bdd_4_lut.init = 16'h0fca;
    LUT4 n23_bdd_3_lut (.A(n23), .B(n34534), .C(tx_byte_index[2]), .Z(n53235)) /* synthesis lut_function=(A (B+(C))+!A !((C)+!B)) */ ;
    defparam n23_bdd_3_lut.init = 16'hacac;
    LUT4 n49411_bdd_3_lut (.A(n49411), .B(tx_word_index[0]), .C(n50860), 
         .Z(n53233)) /* synthesis lut_function=(A ((C)+!B)+!A (B (C))) */ ;
    defparam n49411_bdd_3_lut.init = 16'he2e2;
    LUT4 n52720_bdd_3_lut_41622 (.A(n53869), .B(n52716), .C(tx_word_index[0]), 
         .Z(n53238)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n52720_bdd_3_lut_41622.init = 16'hcaca;
    LUT4 n53239_bdd_3_lut (.A(n53239), .B(n53237), .C(tx_word_index[2]), 
         .Z(n53240)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n53239_bdd_3_lut.init = 16'hcaca;
    LUT4 i1_3_lut_adj_154 (.A(\tx_byte_index[1] ), .B(n34534), .C(n51017), 
         .Z(n3_adj_5116)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i1_3_lut_adj_154.init = 16'hecec;
    FD1S3IX cyc_i_410 (.D(n38167), .CK(sys_clk), .CD(next_state_9__N_4541[6]), 
            .Q(cyc_i)) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=64, LSE_RCOL=6, LSE_LLINE=528, LSE_RLINE=562 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam cyc_i_410.GSR = "ENABLED";
    LUT4 i1_2_lut (.A(\state[5] ), .B(\state[6] ), .Z(n48129)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(366[17:29])
    defparam i1_2_lut.init = 16'heeee;
    LUT4 n25_bdd_4_lut (.A(\VL53L1X_range_mm[4] ), .B(\VL53L1X_range_mm[7] ), 
         .C(\VL53L1X_range_mm[6] ), .D(\VL53L1X_range_mm[5] ), .Z(n53383)) /* synthesis lut_function=(A (C)+!A (B (C (D))+!B (C))) */ ;
    defparam n25_bdd_4_lut.init = 16'hf0b0;
    LUT4 i38914_4_lut (.A(n43332), .B(\tx_byte_index[0] ), .C(\tx_byte_index[1] ), 
         .D(n43302), .Z(n49709)) /* synthesis lut_function=(A (B (C+(D))+!B !(C))+!A (B (C+(D)))) */ ;
    defparam i38914_4_lut.init = 16'hcec2;
    LUT4 i38913_3_lut (.A(n1_adj_5106), .B(n51029), .C(\tx_byte_index[1] ), 
         .Z(n49708)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38913_3_lut.init = 16'hcaca;
    LUT4 n16_bdd_4_lut (.A(n52441), .B(\tx_byte_index[1] ), .C(throttle_val[0]), 
         .D(throttle_val[3]), .Z(n51742)) /* synthesis lut_function=(A (B+!(C (D)+!C !(D)))+!A (B+(C))) */ ;
    defparam n16_bdd_4_lut.init = 16'hdefc;
    PFUMX i31089 (.BLUT(n48537), .ALUT(n71), .C0(\tx_byte_index[0] ), 
          .Z(n6_adj_5117));
    LUT4 i38911_3_lut (.A(n1_adj_5106), .B(n2_adj_5118), .C(\tx_byte_index[1] ), 
         .Z(n49706)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38911_3_lut.init = 16'hcaca;
    LUT4 n11_bdd_4_lut_40642 (.A(throttle_val[4]), .B(throttle_val[5]), 
         .C(throttle_val[7]), .D(throttle_val[6]), .Z(n51743)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A !(B (C)+!B (C (D))))) */ ;
    defparam n11_bdd_4_lut_40642.init = 16'h5a6a;
    LUT4 n50715_bdd_4_lut (.A(\z_linear_velocity[7] ), .B(\z_linear_velocity[4] ), 
         .C(\z_linear_velocity[6] ), .D(\z_linear_velocity[5] ), .Z(n53381)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C)) */ ;
    defparam n50715_bdd_4_lut.init = 16'hf0d0;
    LUT4 n14_bdd_4_lut (.A(n14_adj_5119), .B(\tx_byte_index[1] ), .C(VL53L1X_firm_rdy[0]), 
         .D(VL53L1X_firm_rdy[3]), .Z(n51746)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+!((D)+!C))) */ ;
    defparam n14_bdd_4_lut.init = 16'heefc;
    LUT4 n11_bdd_4_lut_40689 (.A(VL53L1X_firm_rdy[5]), .B(VL53L1X_firm_rdy[4]), 
         .C(VL53L1X_firm_rdy[6]), .D(VL53L1X_firm_rdy[7]), .Z(n51747)) /* synthesis lut_function=(!(A (B (D)+!B !(D))+!A (B (C (D))+!B !(C (D))))) */ ;
    defparam n11_bdd_4_lut_40689.init = 16'h36cc;
    LUT4 i27352_3_lut (.A(\latched_roll[5] ), .B(\latched_roll[7] ), .C(\latched_roll[6] ), 
         .Z(n38035)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i27352_3_lut.init = 16'hc8c8;
    LUT4 n51135_bdd_4_lut (.A(\VL53L1X_range_mm[15] ), .B(\VL53L1X_range_mm[14] ), 
         .C(\VL53L1X_range_mm[13] ), .D(\VL53L1X_range_mm[12] ), .Z(n53396)) /* synthesis lut_function=(A (B (C+(D)))+!A (B)) */ ;
    defparam n51135_bdd_4_lut.init = 16'hccc4;
    LUT4 n52541_bdd_4_lut (.A(\z_linear_velocity[13] ), .B(\z_linear_velocity[15] ), 
         .C(\z_linear_velocity[14] ), .D(\z_linear_velocity[12] ), .Z(n53394)) /* synthesis lut_function=(A (C)+!A (B (C (D))+!B (C))) */ ;
    defparam n52541_bdd_4_lut.init = 16'hf0b0;
    LUT4 tx_byte_index_0__bdd_4_lut_41075 (.A(VL53L1X_chip_id[14]), .B(VL53L1X_chip_id[13]), 
         .C(VL53L1X_chip_id[15]), .D(VL53L1X_chip_id[12]), .Z(n50675)) /* synthesis lut_function=(A (B ((D)+!C)+!B !((D)+!C))+!A (B ((D)+!C))) */ ;
    defparam tx_byte_index_0__bdd_4_lut_41075.init = 16'hcc2c;
    LUT4 i43_4_lut (.A(n20), .B(n27_adj_5120), .C(tx_byte_index[2]), .D(\tx_byte_index[0] ), 
         .Z(n25_c)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(265[13] 275[20])
    defparam i43_4_lut.init = 16'hca0a;
    LUT4 i1_2_lut_adj_155 (.A(state[9]), .B(state[8]), .Z(n44)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(92[29:34])
    defparam i1_2_lut_adj_155.init = 16'h2222;
    LUT4 i27711_4_lut (.A(tx_byte_index[3]), .B(n40), .C(n38267), .D(tx_byte_index[2]), 
         .Z(n38447)) /* synthesis lut_function=(A+(B (C+!(D))+!B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(96[17:30])
    defparam i27711_4_lut.init = 16'hfaee;
    LUT4 i2_3_lut_rep_242_4_lut (.A(state[7]), .B(n52206), .C(state[9]), 
         .D(state[8]), .Z(n52178)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(299[17:22])
    defparam i2_3_lut_rep_242_4_lut.init = 16'hfeff;
    LUT4 i2_4_lut (.A(n49281), .B(n4_adj_5121), .C(n31), .D(n52245), 
         .Z(n7)) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;
    defparam i2_4_lut.init = 16'hccdc;
    LUT4 i1_4_lut_adj_156 (.A(n37479), .B(n52294), .C(n48229), .D(n49106), 
         .Z(n4_adj_5121)) /* synthesis lut_function=(!(A (B+!((D)+!C)))) */ ;
    defparam i1_4_lut_adj_156.init = 16'h7757;
    LUT4 i55_2_lut (.A(state[3]), .B(state[4]), .Z(n31)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;
    defparam i55_2_lut.init = 16'h6666;
    LUT4 i3_4_lut (.A(n52453), .B(n22616), .C(n52454), .D(\state[5] ), 
         .Z(n49106)) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i3_4_lut.init = 16'h0004;
    LUT4 i15445_2_lut (.A(\state[6] ), .B(state[7]), .Z(n22616)) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(218[13] 230[20])
    defparam i15445_2_lut.init = 16'h6666;
    LUT4 n1_bdd_4_lut_41555 (.A(n50864), .B(\tx_byte_index[0] ), .C(\tx_byte_index[1] ), 
         .D(\led_data[4] ), .Z(n53527)) /* synthesis lut_function=(A (B+!(C+!(D)))+!A (B (C)+!B !(C+!(D)))) */ ;
    defparam n1_bdd_4_lut_41555.init = 16'hcbc8;
    LUT4 n2035_bdd_2_lut (.A(n2019[0]), .B(\tx_byte_index[1] ), .Z(n53525)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam n2035_bdd_2_lut.init = 16'h2222;
    LUT4 n53523_bdd_2_lut (.A(n53523), .B(\tx_byte_index[1] ), .Z(n53524)) /* synthesis lut_function=(A+(B)) */ ;
    defparam n53523_bdd_2_lut.init = 16'heeee;
    LUT4 tx_byte_index_1__bdd_4_lut (.A(VL53L1X_chip_id[0]), .B(VL53L1X_chip_id[3]), 
         .C(VL53L1X_chip_id[2]), .D(VL53L1X_chip_id[1]), .Z(n53523)) /* synthesis lut_function=(!(A (B (C+(D)))+!A !(B (C+(D))))) */ ;
    defparam tx_byte_index_1__bdd_4_lut.init = 16'h666a;
    LUT4 n1_bdd_3_lut (.A(n1_adj_5106), .B(n53559), .C(\tx_byte_index[1] ), 
         .Z(n3_adj_5114)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1_bdd_3_lut.init = 16'hcaca;
    LUT4 VL53L1X_chip_id_12__bdd_4_lut (.A(VL53L1X_chip_id[12]), .B(VL53L1X_chip_id[14]), 
         .C(VL53L1X_chip_id[15]), .D(VL53L1X_chip_id[13]), .Z(n53558)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A !(B (C)+!B (C (D))))) */ ;
    defparam VL53L1X_chip_id_12__bdd_4_lut.init = 16'h5a6a;
    LUT4 VL53L1X_chip_id_12__bdd_4_lut_41509 (.A(VL53L1X_chip_id[9]), .B(VL53L1X_chip_id[10]), 
         .C(VL53L1X_chip_id[11]), .D(VL53L1X_chip_id[8]), .Z(n53557)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B !(D)))) */ ;
    defparam VL53L1X_chip_id_12__bdd_4_lut_41509.init = 16'h1fe0;
    LUT4 i2_3_lut_rep_243_4_lut (.A(state[4]), .B(n52208), .C(\state[2] ), 
         .D(state[3]), .Z(n52179)) /* synthesis lut_function=(A+(B+((D)+!C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam i2_3_lut_rep_243_4_lut.init = 16'hffef;
    LUT4 i1_3_lut_adj_157 (.A(\tx_byte_index[1] ), .B(n34534), .C(n50676), 
         .Z(n51)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i1_3_lut_adj_157.init = 16'hecec;
    LUT4 i39285_3_lut (.A(n51), .B(n53874), .C(tx_byte_index[2]), .Z(n9499[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(333[21] 354[28])
    defparam i39285_3_lut.init = 16'hcaca;
    PFUMX i42_adj_158 (.BLUT(n48706), .ALUT(n27_adj_5122), .C0(\tx_byte_index[0] ), 
          .Z(n22_adj_5123));
    LUT4 i39774_2_lut_4_lut (.A(n52184), .B(n47346), .C(n52178), .D(n15182), 
         .Z(n38023)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;
    defparam i39774_2_lut_4_lut.init = 16'h0020;
    LUT4 tx_byte_index_1__bdd_4_lut_40330 (.A(swa_swb_val[5]), .B(swa_swb_val[7]), 
         .C(swa_swb_val[4]), .D(swa_swb_val[6]), .Z(n50975)) /* synthesis lut_function=(A ((C)+!B)+!A !((C+!(D))+!B)) */ ;
    defparam tx_byte_index_1__bdd_4_lut_40330.init = 16'ha6a2;
    LUT4 n11_bdd_4_lut_40316 (.A(swa_swb_val[1]), .B(swa_swb_val[0]), .C(swa_swb_val[3]), 
         .D(swa_swb_val[2]), .Z(n50977)) /* synthesis lut_function=(A (B+!(C))+!A !(B+!(C (D)))) */ ;
    defparam n11_bdd_4_lut_40316.init = 16'h9a8a;
    LUT4 n52718_bdd_4_lut (.A(n52718), .B(\tx_byte_index[1] ), .C(n51353), 
         .D(\tx_byte_index[0] ), .Z(n53869)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam n52718_bdd_4_lut.init = 16'hf0ee;
    LUT4 i1_4_lut_adj_159 (.A(n34729), .B(n52413), .C(n26246), .D(tx_byte_index[2]), 
         .Z(n27740)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(333[21] 354[28])
    defparam i1_4_lut_adj_159.init = 16'hc088;
    LUT4 i1_4_lut_adj_160 (.A(n34729), .B(n47964), .C(n52587), .D(tx_byte_index[2]), 
         .Z(n47966)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_160.init = 16'hc088;
    LUT4 n3_bdd_3_lut (.A(n3_adj_5116), .B(n53870), .C(tx_byte_index[2]), 
         .Z(n53776)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n3_bdd_3_lut.init = 16'hcaca;
    LUT4 i31127_3_lut (.A(n41729), .B(\tx_byte_index[0] ), .C(\tx_byte_index[1] ), 
         .Z(n4)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(96[17:30])
    defparam i31127_3_lut.init = 16'hcaca;
    LUT4 i3_4_lut_adj_161 (.A(n52258), .B(n37731), .C(n23_adj_5124), .D(state[0]), 
         .Z(next_state_9__N_4478[2])) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i3_4_lut_adj_161.init = 16'h0010;
    LUT4 i39809_3_lut_rep_244_4_lut (.A(state[4]), .B(n52208), .C(\state[2] ), 
         .D(state[3]), .Z(n52180)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam i39809_3_lut_rep_244_4_lut.init = 16'h0100;
    PFUMX i40 (.BLUT(n38035), .ALUT(n1406), .C0(\tx_byte_index[0] ), .Z(n21));
    LUT4 i38634_3_lut (.A(n1), .B(n2), .C(\tx_byte_index[1] ), .Z(n49429)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i38634_3_lut.init = 16'hcaca;
    LUT4 i39673_2_lut_rep_237_4_lut_3_lut_4_lut (.A(state[4]), .B(n52208), 
         .C(\state[2] ), .D(state[3]), .Z(n52173)) /* synthesis lut_function=(!(A+(B+(C (D)+!C !(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam i39673_2_lut_rep_237_4_lut_3_lut_4_lut.init = 16'h0110;
    PFUMX i29 (.BLUT(n49483), .ALUT(n49485), .C0(n52375), .Z(n38373));
    LUT4 i1_2_lut_3_lut_4_lut_adj_162 (.A(state[4]), .B(n52451), .C(n52295), 
         .D(n52454), .Z(n27995)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam i1_2_lut_3_lut_4_lut_adj_162.init = 16'hfffe;
    PFUMX i23850 (.BLUT(n48742), .ALUT(n38), .C0(\tx_byte_index[0] ), 
          .Z(n34493));
    LUT4 i1_2_lut_rep_271_3_lut_4_lut (.A(state[4]), .B(n52451), .C(n52295), 
         .D(n48129), .Z(n52207)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam i1_2_lut_rep_271_3_lut_4_lut.init = 16'hfffe;
    LUT4 tx_byte_index_0__bdd_4_lut (.A(\z_linear_velocity[3] ), .B(\z_linear_velocity[2] ), 
         .C(\tx_byte_index[1] ), .D(\z_linear_velocity[1] ), .Z(n53773)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A (C+!(D)))) */ ;
    defparam tx_byte_index_0__bdd_4_lut.init = 16'h0508;
    LUT4 i1_2_lut_rep_270_3_lut_4_lut (.A(state[4]), .B(n52451), .C(n48129), 
         .D(n52454), .Z(n52206)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam i1_2_lut_rep_270_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_272_3_lut_4_lut (.A(state[7]), .B(n52453), .C(n52454), 
         .D(n48129), .Z(n52208)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam i1_2_lut_rep_272_3_lut_4_lut.init = 16'hfffe;
    LUT4 n34481_bdd_4_lut (.A(n34474), .B(\tx_byte_index[1] ), .C(VL53L1X_data_rdy[5]), 
         .D(VL53L1X_data_rdy[6]), .Z(n50859)) /* synthesis lut_function=(A (B+(C))+!A (B+!(C+!(D)))) */ ;
    defparam n34481_bdd_4_lut.init = 16'hedec;
    LUT4 i39904_2_lut_4_lut (.A(state[1]), .B(n52207), .C(state[0]), .D(n37479), 
         .Z(n38167)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)))+!A (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(305[17:25])
    defparam i39904_2_lut_4_lut.init = 16'h02ff;
    LUT4 i27695_4_lut (.A(tx_word_index[4]), .B(n52443), .C(n52398), .D(n25919), 
         .Z(n91)) /* synthesis lut_function=(!(A+(B (C+(D))))) */ ;
    defparam i27695_4_lut.init = 16'h1115;
    LUT4 i1_4_lut_adj_163 (.A(n99_adj_5125), .B(n47964), .C(tx_byte_index[2]), 
         .D(\tx_byte_index[1] ), .Z(n47965)) /* synthesis lut_function=(!(A ((C+!(D))+!B)+!A ((C (D))+!B))) */ ;
    defparam i1_4_lut_adj_163.init = 16'h0c44;
    LUT4 VL53L1X_chip_id_5__bdd_4_lut_41326 (.A(VL53L1X_chip_id[5]), .B(VL53L1X_chip_id[4]), 
         .C(VL53L1X_chip_id[7]), .D(VL53L1X_chip_id[6]), .Z(n51009)) /* synthesis lut_function=(A (B+!(C))+!A !(B+!(C (D)))) */ ;
    defparam VL53L1X_chip_id_5__bdd_4_lut_41326.init = 16'h9a8a;
    PFUMX i38939 (.BLUT(n13_adj_5126), .ALUT(n27_adj_5115), .C0(\tx_byte_index[0] ), 
          .Z(n49734));
    LUT4 z_linear_velocity_13__bdd_4_lut (.A(\z_linear_velocity[13] ), .B(\z_linear_velocity[12] ), 
         .C(\z_linear_velocity[15] ), .D(\z_linear_velocity[14] ), .Z(n51016)) /* synthesis lut_function=(A (B+!(C))+!A !(B+!(C (D)))) */ ;
    defparam z_linear_velocity_13__bdd_4_lut.init = 16'h9a8a;
    LUT4 i1_4_lut_adj_164 (.A(n20), .B(n47964), .C(n6_adj_5117), .D(tx_byte_index[2]), 
         .Z(n47969)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_164.init = 16'hc088;
    LUT4 i1_4_lut_adj_165 (.A(n34534), .B(n47964), .C(n51328), .D(tx_byte_index[2]), 
         .Z(n47967)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_165.init = 16'hc088;
    LUT4 n51351_bdd_3_lut_41189 (.A(n43386), .B(\tx_byte_index[0] ), .C(\tx_byte_index[1] ), 
         .Z(n52715)) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A (B+!(C)))) */ ;
    defparam n51351_bdd_3_lut_41189.init = 16'h3838;
    LUT4 i1_2_lut_adj_166 (.A(VL53L1X_firm_rdy[1]), .B(VL53L1X_firm_rdy[3]), 
         .Z(n48161)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(237[13] 255[20])
    defparam i1_2_lut_adj_166.init = 16'hbbbb;
    PFUMX i38940 (.BLUT(n13_adj_5127), .ALUT(n27_adj_5108), .C0(\tx_byte_index[0] ), 
          .Z(n49735));
    LUT4 i39326_3_lut (.A(n52166), .B(n34665), .C(tx_word_index[0]), .Z(n49376)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(333[21] 354[28])
    defparam i39326_3_lut.init = 16'hcaca;
    PFUMX i40365 (.BLUT(n51327), .ALUT(n51326), .C0(\tx_byte_index[0] ), 
          .Z(n51328));
    PFUMX i38941 (.BLUT(n13_adj_5128), .ALUT(n27_c), .C0(\tx_byte_index[0] ), 
          .Z(n49736));
    LUT4 n51336_bdd_4_lut_41408 (.A(n51336), .B(n51335), .C(\tx_byte_index[0] ), 
         .D(\tx_byte_index[1] ), .Z(n52164)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam n51336_bdd_4_lut_41408.init = 16'hca00;
    PFUMX i40_adj_167 (.BLUT(n37957), .ALUT(n1524[6]), .C0(\tx_byte_index[0] ), 
          .Z(n21_adj_5129));
    LUT4 i41_4_lut (.A(n52434), .B(n304[6]), .C(\tx_byte_index[0] ), .D(tx_word_index[7]), 
         .Z(n18)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(265[13] 275[20])
    defparam i41_4_lut.init = 16'hcac0;
    PFUMX i40362 (.BLUT(n51324), .ALUT(n51323), .C0(n52375), .Z(n51325));
    LUT4 i26515_3_lut (.A(\tx_word_index[1] ), .B(tx_word_index[3]), .C(tx_word_index[2]), 
         .Z(n304[6])) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(237[13] 255[20])
    defparam i26515_3_lut.init = 16'hc8c8;
    LUT4 z_linear_velocity_8__bdd_4_lut_40185 (.A(\z_linear_velocity[8] ), 
         .B(\z_linear_velocity[10] ), .C(\z_linear_velocity[11] ), .D(\z_linear_velocity[9] ), 
         .Z(n51027)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A !(B (C)+!B (C (D))))) */ ;
    defparam z_linear_velocity_8__bdd_4_lut_40185.init = 16'h5a6a;
    LUT4 i38586_4_lut (.A(n52164), .B(n50807), .C(tx_byte_index[2]), .D(n34534), 
         .Z(n49381)) /* synthesis lut_function=(A (B+!(C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;
    defparam i38586_4_lut.init = 16'hcfca;
    LUT4 n51971_bdd_3_lut (.A(n53398), .B(\tx_byte_index[0] ), .C(tx_byte_index[2]), 
         .Z(n51972)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n51971_bdd_3_lut.init = 16'hcaca;
    LUT4 z_linear_velocity_8__bdd_4_lut (.A(\z_linear_velocity[12] ), .B(\z_linear_velocity[14] ), 
         .C(\z_linear_velocity[15] ), .D(\z_linear_velocity[13] ), .Z(n51028)) /* synthesis lut_function=(!(A (B (C)+!B (C (D)))+!A !(B (C)+!B (C (D))))) */ ;
    defparam z_linear_velocity_8__bdd_4_lut.init = 16'h5a6a;
    LUT4 n1_bdd_3_lut_41398 (.A(n1), .B(n53385), .C(tx_byte_index[2]), 
         .Z(n51974)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n1_bdd_3_lut_41398.init = 16'hcaca;
    PFUMX i21 (.BLUT(n50_adj_5130), .ALUT(n5), .C0(\tx_byte_index[0] ), 
          .Z(n7_adj_5131));
    PFUMX i40360 (.BLUT(n51321), .ALUT(n50855), .C0(\tx_byte_index[0] ), 
          .Z(n51322));
    PFUMX i40358 (.BLUT(n51319), .ALUT(n51318), .C0(n52375), .Z(n51320));
    PFUMX i40_adj_168 (.BLUT(n48143), .ALUT(n48199), .C0(\tx_byte_index[0] ), 
          .Z(n38079));
    L6MUX21 i38687 (.D0(n52143), .D1(n52141), .SD(\tx_byte_index[0] ), 
            .Z(n49482));
    PFUMX i41230 (.BLUT(n53075), .ALUT(n25965), .C0(\tx_word_index[1] ), 
          .Z(n53076));
    LUT4 n37942_bdd_4_lut (.A(n37942), .B(n37950), .C(\tx_byte_index[0] ), 
         .D(\tx_byte_index[1] ), .Z(n52165)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (B (C)+!B (C (D)))) */ ;
    defparam n37942_bdd_4_lut.init = 16'hf0ca;
    LUT4 i27721_2_lut (.A(tx_word_index[4]), .B(n38458), .Z(n121)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i27721_2_lut.init = 16'h1111;
    LUT4 n50975_bdd_4_lut_41192 (.A(\latched_roll[6] ), .B(\latched_roll[7] ), 
         .C(\latched_roll[4] ), .D(\latched_roll[5] ), .Z(n52717)) /* synthesis lut_function=(A (B (C (D)+!C !(D))+!B (D))+!A (B (C (D))+!B (D))) */ ;
    defparam n50975_bdd_4_lut_41192.init = 16'hf308;
    LUT4 i1_2_lut_adj_169 (.A(VL53L1X_firm_rdy[5]), .B(VL53L1X_firm_rdy[7]), 
         .Z(n48147)) /* synthesis lut_function=(A+!(B)) */ ;
    defparam i1_2_lut_adj_169.init = 16'hbbbb;
    LUT4 i39293_3_lut_3_lut_then_4_lut (.A(\amc_debug[7] ), .B(\amc_debug[6] ), 
         .C(\amc_debug[5] ), .D(\amc_debug[4] ), .Z(n52496)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)+!C !(D)))+!A !(D))) */ ;
    defparam i39293_3_lut_3_lut_then_4_lut.init = 16'h57a8;
    LUT4 i39293_3_lut_3_lut_else_4_lut (.A(\amc_debug[8] ), .B(n1_adj_5106), 
         .C(\tx_byte_index[1] ), .D(\tx_byte_index[0] ), .Z(n52495)) /* synthesis lut_function=(A (B ((D)+!C)+!B (C (D)))+!A !((C)+!B)) */ ;
    defparam i39293_3_lut_3_lut_else_4_lut.init = 16'hac0c;
    PFUMX i40356 (.BLUT(n48679), .ALUT(n51316), .C0(\tx_byte_index[0] ), 
          .Z(n51317));
    LUT4 i1_2_lut_4_lut_adj_170 (.A(n49426), .B(n49427), .C(tx_word_index[0]), 
         .D(n52414), .Z(n47986)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_2_lut_4_lut_adj_170.init = 16'hca00;
    LUT4 n34679_bdd_4_lut (.A(n48820), .B(n52391), .C(\latched_roll[6] ), 
         .D(\tx_byte_index[0] ), .Z(n52096)) /* synthesis lut_function=(A (B (D)+!B ((D)+!C))+!A !(B+(C+(D)))) */ ;
    defparam n34679_bdd_4_lut.init = 16'haa03;
    CCU2D tx_word_index_6624_add_4_9 (.A0(tx_word_index[7]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43869), .S0(n8[7]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(371[42:62])
    defparam tx_word_index_6624_add_4_9.INIT0 = 16'hfaaa;
    defparam tx_word_index_6624_add_4_9.INIT1 = 16'h0000;
    defparam tx_word_index_6624_add_4_9.INJECT1_0 = "NO";
    defparam tx_word_index_6624_add_4_9.INJECT1_1 = "NO";
    L6MUX21 i38640 (.D0(n21), .D1(n21_adj_5129), .SD(tx_word_index[0]), 
            .Z(n49435));
    CCU2D tx_word_index_6624_add_4_7 (.A0(tx_word_index[5]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(tx_word_index[6]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n43868), .COUT(n43869), .S0(n8[5]), 
          .S1(n8[6]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(371[42:62])
    defparam tx_word_index_6624_add_4_7.INIT0 = 16'hfaaa;
    defparam tx_word_index_6624_add_4_7.INIT1 = 16'hfaaa;
    defparam tx_word_index_6624_add_4_7.INJECT1_0 = "NO";
    defparam tx_word_index_6624_add_4_7.INJECT1_1 = "NO";
    LUT4 i33_3_lut (.A(state[0]), .B(next_state_9__N_4541[6]), .C(state[1]), 
         .Z(n22)) /* synthesis lut_function=(!(A (C)+!A (B+!(C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(218[13] 230[20])
    defparam i33_3_lut.init = 16'h1a1a;
    PFUMX i40042 (.BLUT(n50806), .ALUT(n50805), .C0(\tx_byte_index[0] ), 
          .Z(n50807));
    LUT4 n38079_bdd_3_lut (.A(n38079), .B(n52092), .C(tx_word_index[0]), 
         .Z(n52155)) /* synthesis lut_function=(A (B (C))+!A (B+!(C))) */ ;
    defparam n38079_bdd_3_lut.init = 16'hc5c5;
    LUT4 i1_4_lut_4_lut (.A(\tx_word_index[1] ), .B(\tx_byte_index[0] ), 
         .C(n27), .D(n48692), .Z(n19)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(371[42:62])
    defparam i1_4_lut_4_lut.init = 16'h5140;
    PFUMX mux_4432_Mux_4_i4 (.BLUT(n37943), .ALUT(n37951), .C0(\tx_byte_index[0] ), 
          .Z(n37975));
    LUT4 i1_2_lut_rep_447 (.A(\tx_byte_index[1] ), .B(\tx_byte_index[0] ), 
         .Z(n52383)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(265[13] 275[20])
    defparam i1_2_lut_rep_447.init = 16'h8888;
    LUT4 i33173_3_lut_4_lut (.A(\tx_byte_index[1] ), .B(\tx_byte_index[0] ), 
         .C(tx_byte_index[2]), .D(tx_byte_index[3]), .Z(n9[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(D))+!A !(D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(265[13] 275[20])
    defparam i33173_3_lut_4_lut.init = 16'h7f80;
    LUT4 i33166_2_lut_3_lut (.A(\tx_byte_index[1] ), .B(\tx_byte_index[0] ), 
         .C(tx_byte_index[2]), .Z(n9[2])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(265[13] 275[20])
    defparam i33166_2_lut_3_lut.init = 16'h7878;
    CCU2D tx_word_index_6624_add_4_5 (.A0(tx_word_index[3]), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(tx_word_index[4]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n43867), .COUT(n43868), .S0(n8[3]), 
          .S1(n8[4]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(371[42:62])
    defparam tx_word_index_6624_add_4_5.INIT0 = 16'hfaaa;
    defparam tx_word_index_6624_add_4_5.INIT1 = 16'hfaaa;
    defparam tx_word_index_6624_add_4_5.INJECT1_0 = "NO";
    defparam tx_word_index_6624_add_4_5.INJECT1_1 = "NO";
    LUT4 i27273_3_lut_4_lut (.A(VL53L1X_chip_id[1]), .B(VL53L1X_chip_id[3]), 
         .C(VL53L1X_chip_id[2]), .D(VL53L1X_chip_id[0]), .Z(n37950)) /* synthesis lut_function=(A (C)+!A (B (C (D))+!B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(237[13] 255[20])
    defparam i27273_3_lut_4_lut.init = 16'hf0b0;
    FD1S3IX state_i9 (.D(next_state_9__N_4478[9]), .CK(sys_clk), .CD(resetn_derived_2), 
            .Q(state[9])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=64, LSE_RCOL=6, LSE_LLINE=528, LSE_RLINE=562 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam state_i9.GSR = "ENABLED";
    LUT4 n42194_bdd_4_lut (.A(\VL53L1X_range_mm[12] ), .B(\VL53L1X_range_mm[15] ), 
         .C(\VL53L1X_range_mm[13] ), .D(\VL53L1X_range_mm[14] ), .Z(n51336)) /* synthesis lut_function=(A (C)+!A !(B (C+!(D))+!B !(C))) */ ;
    defparam n42194_bdd_4_lut.init = 16'hb4b0;
    FD1S3IX state_i8 (.D(next_state_9__N_4478[8]), .CK(sys_clk), .CD(resetn_derived_2), 
            .Q(state[8])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=64, LSE_RCOL=6, LSE_LLINE=528, LSE_RLINE=562 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam state_i8.GSR = "ENABLED";
    FD1S3IX state_i7 (.D(next_state_9__N_4478[7]), .CK(sys_clk), .CD(resetn_derived_2), 
            .Q(state[7])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=64, LSE_RCOL=6, LSE_LLINE=528, LSE_RLINE=562 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam state_i7.GSR = "ENABLED";
    FD1S3IX state_i6 (.D(next_state_9__N_4478[6]), .CK(sys_clk), .CD(resetn_derived_2), 
            .Q(\state[6] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=64, LSE_RCOL=6, LSE_LLINE=528, LSE_RLINE=562 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam state_i6.GSR = "ENABLED";
    FD1S3IX state_i5 (.D(next_state_9__N_4478[5]), .CK(sys_clk), .CD(resetn_derived_2), 
            .Q(\state[5] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=64, LSE_RCOL=6, LSE_LLINE=528, LSE_RLINE=562 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam state_i5.GSR = "ENABLED";
    FD1S3IX state_i4 (.D(next_state_9__N_4478[4]), .CK(sys_clk), .CD(resetn_derived_2), 
            .Q(state[4])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=64, LSE_RCOL=6, LSE_LLINE=528, LSE_RLINE=562 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam state_i4.GSR = "ENABLED";
    FD1S3IX state_i3 (.D(next_state_9__N_4478[3]), .CK(sys_clk), .CD(resetn_derived_2), 
            .Q(state[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=64, LSE_RCOL=6, LSE_LLINE=528, LSE_RLINE=562 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam state_i3.GSR = "ENABLED";
    FD1S3IX state_i2 (.D(next_state_9__N_4478[2]), .CK(sys_clk), .CD(resetn_derived_2), 
            .Q(\state[2] )) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=64, LSE_RCOL=6, LSE_LLINE=528, LSE_RLINE=562 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam state_i2.GSR = "ENABLED";
    FD1S3IX state_i1 (.D(next_state_9__N_4478[1]), .CK(sys_clk), .CD(resetn_derived_2), 
            .Q(state[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=64, LSE_RCOL=6, LSE_LLINE=528, LSE_RLINE=562 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam state_i1.GSR = "ENABLED";
    FD1S3AX adr_i_i3 (.D(n52180), .CK(sys_clk), .Q(adr_i[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=64, LSE_RCOL=6, LSE_LLINE=528, LSE_RLINE=562 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam adr_i_i3.GSR = "ENABLED";
    FD1S3AX adr_i_i2 (.D(n52173), .CK(sys_clk), .Q(adr_i[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=64, LSE_RCOL=6, LSE_LLINE=528, LSE_RLINE=562 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam adr_i_i2.GSR = "ENABLED";
    FD1P3AX dat_i_i5 (.D(next_dat_i_15__N_4452[4]), .SP(sys_clk_enable_246), 
            .CK(sys_clk), .Q(dat_i[5])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=64, LSE_RCOL=6, LSE_LLINE=528, LSE_RLINE=562 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam dat_i_i5.GSR = "ENABLED";
    LUT4 i39746_2_lut (.A(tx_word_index[3]), .B(\tx_word_index[1] ), .Z(n49682)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(333[21] 354[28])
    defparam i39746_2_lut.init = 16'hbbbb;
    LUT4 n48141_bdd_3_lut_40331_4_lut (.A(swa_swb_val[5]), .B(swa_swb_val[7]), 
         .C(swa_swb_val[6]), .D(swa_swb_val[4]), .Z(n51271)) /* synthesis lut_function=(A (C)+!A (B (C (D))+!B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(237[13] 255[20])
    defparam n48141_bdd_3_lut_40331_4_lut.init = 16'hf0b0;
    LUT4 i1_2_lut_3_lut_adj_171 (.A(swa_swb_val[5]), .B(swa_swb_val[7]), 
         .C(swa_swb_val[6]), .Z(n48143)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(237[13] 255[20])
    defparam i1_2_lut_3_lut_adj_171.init = 16'hfbfb;
    LUT4 i1_2_lut_rep_455 (.A(\latched_roll[5] ), .B(\latched_roll[7] ), 
         .Z(n52391)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(237[13] 255[20])
    defparam i1_2_lut_rep_455.init = 16'hbbbb;
    LUT4 n48141_bdd_3_lut_4_lut (.A(\latched_roll[5] ), .B(\latched_roll[7] ), 
         .C(\latched_roll[6] ), .D(\latched_roll[4] ), .Z(n51272)) /* synthesis lut_function=(A (C)+!A (B (C (D))+!B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(237[13] 255[20])
    defparam n48141_bdd_3_lut_4_lut.init = 16'hf0b0;
    LUT4 i39297_3_lut_3_lut (.A(tx_word_index[0]), .B(n25_c), .C(n52165), 
         .Z(n49431)) /* synthesis lut_function=(A (C)+!A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(371[42:62])
    defparam i39297_3_lut_3_lut.init = 16'he4e4;
    LUT4 i31055_1_lut_rep_459 (.A(\tx_byte_index[0] ), .Z(n52395)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam i31055_1_lut_rep_459.init = 16'h5555;
    LUT4 n314_bdd_4_lut (.A(n304[6]), .B(tx_word_index[0]), .C(n50907), 
         .D(\tx_byte_index[0] ), .Z(n1_adj_5106)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(C+(D)))+!A !(B (C+(D))+!B !((D)+!C)))) */ ;
    defparam n314_bdd_4_lut.init = 16'h66f0;
    LUT4 i2_3_lut_4_lut_4_lut_4_lut (.A(\tx_byte_index[0] ), .B(\led_data[1] ), 
         .C(\led_data[2] ), .D(\led_data[3] ), .Z(n48861)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam i2_3_lut_4_lut_4_lut_4_lut.init = 16'hfdff;
    CCU2D tx_word_index_6624_add_4_3 (.A0(\tx_word_index[1] ), .B0(GND_net), 
          .C0(GND_net), .D0(GND_net), .A1(tx_word_index[2]), .B1(GND_net), 
          .C1(GND_net), .D1(GND_net), .CIN(n43866), .COUT(n43867), .S0(n8[1]), 
          .S1(n8[2]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(371[42:62])
    defparam tx_word_index_6624_add_4_3.INIT0 = 16'hfaaa;
    defparam tx_word_index_6624_add_4_3.INIT1 = 16'hfaaa;
    defparam tx_word_index_6624_add_4_3.INJECT1_0 = "NO";
    defparam tx_word_index_6624_add_4_3.INJECT1_1 = "NO";
    PFUMX i31617 (.BLUT(n42210), .ALUT(n42214), .C0(\tx_byte_index[0] ), 
          .Z(n2_adj_5118));
    LUT4 i26369_2_lut_rep_462 (.A(tx_byte_index[3]), .B(\tx_byte_index[1] ), 
         .Z(n52398)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i26369_2_lut_rep_462.init = 16'heeee;
    LUT4 i2_3_lut_3_lut_3_lut_4_lut (.A(tx_byte_index[3]), .B(\tx_byte_index[1] ), 
         .C(n25919), .D(tx_word_index[4]), .Z(n48839)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;
    defparam i2_3_lut_3_lut_3_lut_4_lut.init = 16'h0010;
    CCU2D tx_word_index_6624_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(tx_word_index[0]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n43866), .S1(n8[0]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(371[42:62])
    defparam tx_word_index_6624_add_4_1.INIT0 = 16'hF000;
    defparam tx_word_index_6624_add_4_1.INIT1 = 16'h0555;
    defparam tx_word_index_6624_add_4_1.INJECT1_0 = "NO";
    defparam tx_word_index_6624_add_4_1.INJECT1_1 = "NO";
    LUT4 i38806_2_lut_rep_463 (.A(\tx_byte_index[1] ), .B(\tx_byte_index[0] ), 
         .Z(n52399)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(265[13] 275[20])
    defparam i38806_2_lut_rep_463.init = 16'h2222;
    LUT4 n43221_bdd_4_lut (.A(n43221), .B(n43225), .C(\tx_byte_index[0] ), 
         .D(\tx_byte_index[1] ), .Z(n52167)) /* synthesis lut_function=(A (B (C+!(D))+!B (C (D)+!C !(D)))+!A (B (C)+!B (C (D)))) */ ;
    defparam n43221_bdd_4_lut.init = 16'hf0ca;
    LUT4 i39696_2_lut_rep_336_3_lut (.A(\tx_byte_index[1] ), .B(\tx_byte_index[0] ), 
         .C(tx_byte_index[2]), .Z(n52272)) /* synthesis lut_function=(!(A (C)+!A (B (C)))) */ ;
    defparam i39696_2_lut_rep_336_3_lut.init = 16'h1f1f;
    LUT4 i26036_2_lut (.A(swa_swb_val[0]), .B(swa_swb_val[1]), .Z(n10)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(237[13] 255[20])
    defparam i26036_2_lut.init = 16'h8888;
    LUT4 i22237_1_lut_rep_442 (.A(tx_word_index[2]), .Z(n52378)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(371[42:62])
    defparam i22237_1_lut_rep_442.init = 16'h5555;
    LUT4 i1_2_lut_3_lut_adj_172 (.A(\VL53L1X_range_mm[13] ), .B(\VL53L1X_range_mm[14] ), 
         .C(\VL53L1X_range_mm[15] ), .Z(n50_adj_5130)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;
    defparam i1_2_lut_3_lut_adj_172.init = 16'he0e0;
    PFUMX i40021 (.BLUT(n50747), .ALUT(n50746), .C0(\tx_byte_index[0] ), 
          .Z(n1));
    LUT4 n48198_bdd_4_lut (.A(n52359), .B(swa_swb_val[3]), .C(n50884), 
         .D(\tx_byte_index[0] ), .Z(n52160)) /* synthesis lut_function=(A (B (C+(D))+!B !((D)+!C))+!A !((D)+!C)) */ ;
    defparam n48198_bdd_4_lut.init = 16'h88f0;
    LUT4 i2_3_lut (.A(tx_word_index[4]), .B(tx_byte_index[3]), .C(tx_word_index[0]), 
         .Z(n47964)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(371[42:62])
    defparam i2_3_lut.init = 16'h0202;
    LUT4 i39692_2_lut (.A(tx_byte_index[2]), .B(\tx_byte_index[0] ), .Z(n49697)) /* synthesis lut_function=(!(A (B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(333[21] 354[28])
    defparam i39692_2_lut.init = 16'h7777;
    LUT4 i15480_4_lut (.A(n22_adj_5123), .B(n34493), .C(tx_word_index[0]), 
         .D(n52383), .Z(n25954)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(333[21] 354[28])
    defparam i15480_4_lut.init = 16'hfaca;
    LUT4 i106_3_lut (.A(n18), .B(n49), .C(tx_byte_index[2]), .Z(n99_adj_5125)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam i106_3_lut.init = 16'hcaca;
    LUT4 i39758_2_lut_rep_471 (.A(tx_word_index[2]), .B(\tx_word_index[1] ), 
         .Z(n52407)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(333[21] 354[28])
    defparam i39758_2_lut_rep_471.init = 16'hdddd;
    LUT4 i32_3_lut_4_lut (.A(\amc_debug[2] ), .B(\amc_debug[1] ), .C(\amc_debug[3] ), 
         .D(\amc_debug[0] ), .Z(n41729)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B !(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(184[18:27])
    defparam i32_3_lut_4_lut.init = 16'h1fe0;
    LUT4 i1_2_lut_3_lut_adj_173 (.A(\amc_debug[2] ), .B(\amc_debug[1] ), 
         .C(\amc_debug[3] ), .Z(n89)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(184[18:27])
    defparam i1_2_lut_3_lut_adj_173.init = 16'he0e0;
    LUT4 n43309_bdd_4_lut (.A(n43309), .B(\tx_byte_index[1] ), .C(n53773), 
         .D(\tx_byte_index[0] ), .Z(n53870)) /* synthesis lut_function=(A (C+!(D))+!A (B (C+!(D))+!B (C (D)))) */ ;
    defparam n43309_bdd_4_lut.init = 16'hf0ee;
    LUT4 i1_4_lut_adj_174 (.A(n50956), .B(n48081), .C(n27651), .D(n30), 
         .Z(next_dat_i_15__N_4452[4])) /* synthesis lut_function=(A (B (C))+!A (B (C+!(D)))) */ ;
    defparam i1_4_lut_adj_174.init = 16'hc0c4;
    LUT4 i1_2_lut_3_lut_adj_175 (.A(\amc_debug[5] ), .B(\amc_debug[6] ), 
         .C(\amc_debug[7] ), .Z(n65)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(184[18:27])
    defparam i1_2_lut_3_lut_adj_175.init = 16'he0e0;
    LUT4 i15764_2_lut (.A(\tx_byte_index[1] ), .B(n51047), .Z(n26246)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(333[21] 354[28])
    defparam i15764_2_lut.init = 16'hbbbb;
    PFUMX i24133 (.BLUT(n48828), .ALUT(n49185), .C0(\tx_byte_index[0] ), 
          .Z(n23_adj_5139));
    LUT4 n11_bdd_4_lut_40002 (.A(n52456), .B(\tx_byte_index[1] ), .C(yaw_val[0]), 
         .D(yaw_val[3]), .Z(n50718)) /* synthesis lut_function=(A (B+!(C (D)+!C !(D)))+!A (B+(C))) */ ;
    defparam n11_bdd_4_lut_40002.init = 16'hdefc;
    LUT4 n11_bdd_4_lut_40019 (.A(yaw_val[4]), .B(yaw_val[7]), .C(yaw_val[6]), 
         .D(yaw_val[5]), .Z(n50719)) /* synthesis lut_function=(!(A (B (C+(D)))+!A !(B (C+(D))))) */ ;
    defparam n11_bdd_4_lut_40019.init = 16'h666a;
    PFUMX i40924 (.BLUT(n52495), .ALUT(n52496), .C0(tx_byte_index[2]), 
          .Z(n52497));
    LUT4 i39317_3_lut_4_lut (.A(tx_word_index[0]), .B(tx_byte_index[2]), 
         .C(n49431), .D(n49429), .Z(n5_adj_5140)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;
    defparam i39317_3_lut_4_lut.init = 16'hf2d0;
    LUT4 i25875_4_lut_4_lut (.A(tx_byte_index[3]), .B(tx_byte_index[2]), 
         .C(n6_adj_5141), .D(n40), .Z(n9354[6])) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam i25875_4_lut_4_lut.init = 16'h5140;
    LUT4 i2_3_lut_3_lut_3_lut (.A(tx_byte_index[3]), .B(n53078), .C(tx_word_index[4]), 
         .Z(n49085)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam i2_3_lut_3_lut_3_lut.init = 16'h0404;
    LUT4 i39830_2_lut_rep_477 (.A(tx_byte_index[3]), .B(tx_word_index[4]), 
         .Z(n52413)) /* synthesis lut_function=(!(A+(B))) */ ;
    defparam i39830_2_lut_rep_477.init = 16'h1111;
    LUT4 i1_2_lut_3_lut_adj_176 (.A(tx_byte_index[3]), .B(tx_word_index[4]), 
         .C(n51320), .Z(n27742)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_176.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_177 (.A(tx_byte_index[3]), .B(tx_word_index[4]), 
         .C(n51325), .Z(n27743)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_177.init = 16'h1010;
    LUT4 i1_2_lut_3_lut_adj_178 (.A(tx_byte_index[3]), .B(tx_word_index[4]), 
         .C(n25959), .Z(n27741)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i1_2_lut_3_lut_adj_178.init = 16'h1010;
    LUT4 i2_2_lut_3_lut (.A(tx_byte_index[3]), .B(tx_word_index[4]), .C(n51631), 
         .Z(n48972)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i2_2_lut_3_lut.init = 16'h1010;
    LUT4 i2_2_lut_3_lut_adj_179 (.A(tx_byte_index[3]), .B(tx_word_index[4]), 
         .C(n48486), .Z(n48928)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i2_2_lut_3_lut_adj_179.init = 16'h1010;
    LUT4 i2_2_lut_3_lut_adj_180 (.A(tx_byte_index[3]), .B(tx_word_index[4]), 
         .C(n53240), .Z(n48969)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;
    defparam i2_2_lut_3_lut_adj_180.init = 16'h1010;
    LUT4 i2_3_lut_rep_478 (.A(tx_word_index[4]), .B(tx_byte_index[3]), .C(tx_word_index[2]), 
         .Z(n52414)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(371[42:62])
    defparam i2_3_lut_rep_478.init = 16'h0202;
    LUT4 i1_2_lut_4_lut_adj_181 (.A(tx_word_index[4]), .B(tx_byte_index[3]), 
         .C(tx_word_index[2]), .D(n49401), .Z(n47988)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(371[42:62])
    defparam i1_2_lut_4_lut_adj_181.init = 16'h0200;
    LUT4 i1_2_lut_4_lut_adj_182 (.A(tx_word_index[4]), .B(tx_byte_index[3]), 
         .C(tx_word_index[2]), .D(n51975), .Z(n47990)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(371[42:62])
    defparam i1_2_lut_4_lut_adj_182.init = 16'h0200;
    LUT4 i1_2_lut_4_lut_adj_183 (.A(tx_word_index[4]), .B(tx_byte_index[3]), 
         .C(tx_word_index[2]), .D(n49712), .Z(n47989)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(371[42:62])
    defparam i1_2_lut_4_lut_adj_183.init = 16'h0200;
    LUT4 i1_2_lut_3_lut_adj_184 (.A(\z_linear_velocity[9] ), .B(\z_linear_velocity[10] ), 
         .C(\z_linear_velocity[11] ), .Z(n6)) /* synthesis lut_function=(!(A+(B+!(C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(237[13] 255[20])
    defparam i1_2_lut_3_lut_adj_184.init = 16'h1010;
    LUT4 i26986_2_lut_3_lut (.A(\z_linear_velocity[13] ), .B(\z_linear_velocity[15] ), 
         .C(\z_linear_velocity[14] ), .Z(n1_adj_5113)) /* synthesis lut_function=(!(A+((C)+!B))) */ ;
    defparam i26986_2_lut_3_lut.init = 16'h0404;
    LUT4 i39_4_lut (.A(n18), .B(\led_data[3] ), .C(tx_byte_index[2]), 
         .D(n4_adj_5142), .Z(n24)) /* synthesis lut_function=(A (B ((D)+!C)+!B !(C))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(265[13] 275[20])
    defparam i39_4_lut.init = 16'hca0a;
    LUT4 i1_3_lut_adj_185 (.A(\tx_byte_index[0] ), .B(\led_data[1] ), .C(\led_data[2] ), 
         .Z(n4_adj_5142)) /* synthesis lut_function=(A (B+(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(265[13] 275[20])
    defparam i1_3_lut_adj_185.init = 16'ha8a8;
    LUT4 i40_3_lut (.A(n18), .B(n52563), .C(\tx_byte_index[1] ), .Z(n40)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(96[17:30])
    defparam i40_3_lut.init = 16'hcaca;
    LUT4 i27564_2_lut (.A(n37975), .B(\tx_byte_index[1] ), .Z(n38267)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i27564_2_lut.init = 16'heeee;
    LUT4 i1_4_lut_adj_186 (.A(\tx_byte_index[1] ), .B(\led_data[0] ), .C(\led_data[2] ), 
         .D(n52267), .Z(n27_adj_5120)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(265[13] 275[20])
    defparam i1_4_lut_adj_186.init = 16'hfaea;
    LUT4 i31612_4_lut_4_lut (.A(\VL53L1X_range_mm[12] ), .B(\VL53L1X_range_mm[13] ), 
         .C(\VL53L1X_range_mm[14] ), .D(\VL53L1X_range_mm[15] ), .Z(n42210)) /* synthesis lut_function=(!(A (B (D)+!B (C (D)))+!A !(B (D)+!B (C (D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(155[9:25])
    defparam i31612_4_lut_4_lut.init = 16'h56aa;
    LUT4 i1_2_lut_rep_392 (.A(latched_pitch[5]), .B(latched_pitch[7]), .Z(n52328)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(237[13] 255[20])
    defparam i1_2_lut_rep_392.init = 16'hbbbb;
    LUT4 mux_285_Mux_0_i14_3_lut (.A(VL53L1X_firm_rdy[0]), .B(VL53L1X_firm_rdy[2]), 
         .C(VL53L1X_firm_rdy[1]), .Z(n14_adj_5119)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(237[13] 255[20])
    defparam mux_285_Mux_0_i14_3_lut.init = 16'h5656;
    LUT4 swa_swb_val_1__bdd_3_lut (.A(swa_swb_val[1]), .B(swa_swb_val[2]), 
         .C(swa_swb_val[0]), .Z(n51157)) /* synthesis lut_function=(!(A (C)+!A (B (C)+!B !(C)))) */ ;
    defparam swa_swb_val_1__bdd_3_lut.init = 16'h1e1e;
    LUT4 i1_3_lut_adj_187 (.A(\tx_byte_index[1] ), .B(n34729), .C(n23_adj_5139), 
         .Z(n3)) /* synthesis lut_function=(A (B+(C))+!A (B)) */ ;
    defparam i1_3_lut_adj_187.init = 16'hecec;
    LUT4 i1_2_lut_3_lut_adj_188 (.A(VL53L1X_data_rdy[1]), .B(VL53L1X_data_rdy[2]), 
         .C(VL53L1X_data_rdy[3]), .Z(n11)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(161[9:25])
    defparam i1_2_lut_3_lut_adj_188.init = 16'he0e0;
    LUT4 i23_3_lut_4_lut (.A(VL53L1X_data_rdy[1]), .B(VL53L1X_data_rdy[2]), 
         .C(VL53L1X_data_rdy[3]), .D(VL53L1X_data_rdy[0]), .Z(n34503)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B !(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(161[9:25])
    defparam i23_3_lut_4_lut.init = 16'h1fe0;
    LUT4 i1_2_lut_rep_483 (.A(VL53L1X_data_rdy[5]), .B(VL53L1X_data_rdy[6]), 
         .Z(n52419)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(161[9:25])
    defparam i1_2_lut_rep_483.init = 16'heeee;
    LUT4 i1_2_lut_3_lut_adj_189 (.A(VL53L1X_data_rdy[5]), .B(VL53L1X_data_rdy[6]), 
         .C(VL53L1X_data_rdy[7]), .Z(n3_adj_5112)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(161[9:25])
    defparam i1_2_lut_3_lut_adj_189.init = 16'he0e0;
    LUT4 i27266_3_lut_4_lut (.A(VL53L1X_chip_id[5]), .B(VL53L1X_chip_id[7]), 
         .C(VL53L1X_chip_id[6]), .D(VL53L1X_chip_id[4]), .Z(n37942)) /* synthesis lut_function=(A (C)+!A (B (C (D))+!B (C))) */ ;
    defparam i27266_3_lut_4_lut.init = 16'hf0b0;
    PFUMX i40003 (.BLUT(n50720), .ALUT(n50718), .C0(\tx_byte_index[0] ), 
          .Z(n50721));
    LUT4 THRE_I_0_1_lut (.A(next_state_9__N_4551[6]), .Z(txrdy_n_c_7)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_core.v(320[23:28])
    defparam THRE_I_0_1_lut.init = 16'h5555;
    LUT4 i34_4_lut_3_lut (.A(state[1]), .B(next_state_9__N_4541[6]), .C(\state[2] ), 
         .Z(n23_adj_5124)) /* synthesis lut_function=(!(A ((C)+!B)+!A (B+!(C)))) */ ;
    defparam i34_4_lut_3_lut.init = 16'h1818;
    LUT4 i1_2_lut_4_lut_adj_190 (.A(n49381), .B(n53776), .C(tx_word_index[0]), 
         .D(n52414), .Z(n47985)) /* synthesis lut_function=(A (B (D)+!B !(C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_2_lut_4_lut_adj_190.init = 16'hca00;
    LUT4 i20_3_lut (.A(n18), .B(n7_adj_5131), .C(\tx_byte_index[1] ), 
         .Z(n38325)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(96[17:30])
    defparam i20_3_lut.init = 16'hcaca;
    LUT4 mux_4456_Mux_5_i3_3_lut (.A(n18), .B(n52599), .C(\tx_byte_index[1] ), 
         .Z(n38329)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(265[13] 275[20])
    defparam mux_4456_Mux_5_i3_3_lut.init = 16'hcaca;
    LUT4 i39806_4_lut (.A(n47346), .B(n52184), .C(n44893), .D(n52180), 
         .Z(sys_clk_enable_236)) /* synthesis lut_function=(!(A (B)+!A (B (C+(D))))) */ ;
    defparam i39806_4_lut.init = 16'h3337;
    LUT4 i33159_2_lut (.A(\tx_byte_index[1] ), .B(\tx_byte_index[0] ), .Z(n9[1])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam i33159_2_lut.init = 16'h6666;
    LUT4 i2_3_lut_rep_405 (.A(\state[6] ), .B(state[7]), .C(state[4]), 
         .Z(n52341)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i2_3_lut_rep_405.init = 16'hfefe;
    LUT4 i1_2_lut_rep_322_4_lut (.A(\state[6] ), .B(state[7]), .C(state[4]), 
         .D(\state[5] ), .Z(n52258)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i1_2_lut_rep_322_4_lut.init = 16'hfffe;
    LUT4 i25974_2_lut_rep_406 (.A(state[1]), .B(state[0]), .Z(n52342)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i25974_2_lut_rep_406.init = 16'heeee;
    LUT4 tx_word_index_3__bdd_4_lut_40020 (.A(tx_word_index[3]), .B(tx_word_index[0]), 
         .C(tx_word_index[2]), .D(\tx_word_index[1] ), .Z(n50746)) /* synthesis lut_function=(A (B (C)+!B (C (D)))+!A (C)) */ ;
    defparam tx_word_index_3__bdd_4_lut_40020.init = 16'hf0d0;
    LUT4 i27471_2_lut_3_lut_4_lut (.A(state[1]), .B(state[0]), .C(n52451), 
         .D(n52453), .Z(n38171)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i27471_2_lut_3_lut_4_lut.init = 16'hfffe;
    LUT4 mux_188_Mux_0_i14_3_lut (.A(\latched_roll[4] ), .B(\latched_roll[6] ), 
         .C(\latched_roll[5] ), .Z(n14_adj_5144)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(237[13] 255[20])
    defparam mux_188_Mux_0_i14_3_lut.init = 16'h5656;
    LUT4 i37558_2_lut_rep_321_3_lut (.A(state[1]), .B(state[0]), .C(state[9]), 
         .Z(n52257)) /* synthesis lut_function=(A+(B+(C))) */ ;
    defparam i37558_2_lut_rep_321_3_lut.init = 16'hfefe;
    LUT4 mux_204_Mux_0_i14_3_lut (.A(latched_pitch[4]), .B(latched_pitch[6]), 
         .C(latched_pitch[5]), .Z(n14_adj_5145)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(237[13] 255[20])
    defparam mux_204_Mux_0_i14_3_lut.init = 16'h5656;
    LUT4 mux_205_Mux_0_i14_3_lut (.A(latched_pitch[0]), .B(latched_pitch[2]), 
         .C(latched_pitch[1]), .Z(n14)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(237[13] 255[20])
    defparam mux_205_Mux_0_i14_3_lut.init = 16'h5656;
    LUT4 mux_220_Mux_0_i14_3_lut (.A(swa_swb_val[4]), .B(swa_swb_val[6]), 
         .C(swa_swb_val[5]), .Z(n14_adj_5146)) /* synthesis lut_function=(!(A (B+(C))+!A !(B+(C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(237[13] 255[20])
    defparam mux_220_Mux_0_i14_3_lut.init = 16'h5656;
    LUT4 i1_2_lut_4_lut_adj_191 (.A(n49423), .B(n49424), .C(tx_word_index[0]), 
         .D(n52414), .Z(n47987)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+!(D))+!B !(D)))) */ ;
    defparam i1_2_lut_4_lut_adj_191.init = 16'h3500;
    LUT4 tx_word_index_3__bdd_4_lut_40528 (.A(tx_word_index[4]), .B(tx_word_index[6]), 
         .C(tx_word_index[5]), .D(tx_word_index[7]), .Z(n50747)) /* synthesis lut_function=(A (B)+!A (B (C+!(D)))) */ ;
    defparam tx_word_index_3__bdd_4_lut_40528.init = 16'hc8cc;
    LUT4 i1_2_lut_rep_486 (.A(yaw_val[5]), .B(yaw_val[7]), .Z(n52422)) /* synthesis lut_function=(A+!(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(237[13] 255[20])
    defparam i1_2_lut_rep_486.init = 16'hbbbb;
    LUT4 yaw_val_3__bdd_2_lut_3_lut (.A(yaw_val[5]), .B(yaw_val[7]), .C(yaw_val[6]), 
         .Z(n51042)) /* synthesis lut_function=(A+((C)+!B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(237[13] 255[20])
    defparam yaw_val_3__bdd_2_lut_3_lut.init = 16'hfbfb;
    LUT4 i1_2_lut_4_lut_adj_192 (.A(n52451), .B(n52208), .C(state[4]), 
         .D(n7), .Z(n40166)) /* synthesis lut_function=(!(A (D)+!A (B (D)+!B (C+(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam i1_2_lut_4_lut_adj_192.init = 16'h00ef;
    LUT4 i2_4_lut_adj_193 (.A(n52255), .B(n52179), .C(n123_c), .D(n86), 
         .Z(n48589)) /* synthesis lut_function=(A ((D)+!B)+!A ((C+(D))+!B)) */ ;
    defparam i2_4_lut_adj_193.init = 16'hff73;
    LUT4 i1_4_lut_adj_194 (.A(n34534), .B(n81), .C(n52399), .D(tx_byte_index[2]), 
         .Z(n86)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_194.init = 16'hc088;
    LUT4 i1_4_lut_adj_195 (.A(n85), .B(n48081), .C(n52255), .D(n37), 
         .Z(next_dat_i_15__N_4452[2])) /* synthesis lut_function=(A (B)+!A !((C+!(D))+!B)) */ ;
    defparam i1_4_lut_adj_195.init = 16'h8c88;
    LUT4 i1_4_lut_adj_196 (.A(n20), .B(n81), .C(n52383), .D(tx_byte_index[2]), 
         .Z(n85)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;
    defparam i1_4_lut_adj_196.init = 16'hc088;
    LUT4 i1_4_lut_adj_197 (.A(n34729), .B(n81), .C(\tx_byte_index[1] ), 
         .D(tx_byte_index[2]), .Z(n27734)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(226[60:96])
    defparam i1_4_lut_adj_197.init = 16'hc088;
    LUT4 i1_4_lut_adj_198 (.A(n49126), .B(n48081), .C(n52255), .D(n39_adj_5147), 
         .Z(next_dat_i_15__N_4452[6])) /* synthesis lut_function=(A (B)+!A !((C+!(D))+!B)) */ ;
    defparam i1_4_lut_adj_198.init = 16'h8c88;
    LUT4 i36_4_lut_4_lut (.A(next_state_9__N_4571[5]), .B(state[3]), .C(next_state_9__N_4531[5]), 
         .D(state[8]), .Z(n20_adj_5148)) /* synthesis lut_function=(!(A (B ((D)+!C)+!B !(D))+!A (((D)+!C)+!B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(218[13] 230[20])
    defparam i36_4_lut_4_lut.init = 16'h22c0;
    LUT4 i13_3_lut_4_lut (.A(\VL53L1X_range_mm[9] ), .B(\VL53L1X_range_mm[10] ), 
         .C(\VL53L1X_range_mm[11] ), .D(\VL53L1X_range_mm[8] ), .Z(n42214)) /* synthesis lut_function=(!(A (C (D)+!C !(D))+!A (B (C (D)+!C !(D))+!B !(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(155[9:25])
    defparam i13_3_lut_4_lut.init = 16'h1fe0;
    PFUMX i41038 (.BLUT(n52717), .ALUT(n50975), .C0(\tx_word_index[1] ), 
          .Z(n52718));
    L6MUX21 i40200 (.D0(n51046), .D1(n51043), .SD(tx_word_index[0]), .Z(n51047));
    PFUMX i40198 (.BLUT(n51045), .ALUT(n51044), .C0(\tx_byte_index[0] ), 
          .Z(n51046));
    L6MUX21 i40871 (.D0(n52097), .D1(n52155), .SD(\tx_word_index[1] ), 
            .Z(n26269));
    L6MUX21 i25101 (.D0(n108), .D1(n117), .SD(n49682), .Z(n41_adj_5149));
    PFUMX i40869 (.BLUT(n52096), .ALUT(n52095), .C0(tx_word_index[0]), 
          .Z(n52097));
    L6MUX21 i169 (.D0(n108_adj_5150), .D1(n117_adj_5151), .SD(n49682), 
            .Z(n123_c));
    LUT4 i27274_3_lut (.A(VL53L1X_chip_id[1]), .B(VL53L1X_chip_id[3]), .C(VL53L1X_chip_id[2]), 
         .Z(n37951)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i27274_3_lut.init = 16'hc8c8;
    PFUMX i167 (.BLUT(n47985), .ALUT(n48969), .C0(tx_word_index[3]), .Z(n117_adj_5151));
    LUT4 i27267_3_lut (.A(VL53L1X_chip_id[5]), .B(VL53L1X_chip_id[7]), .C(VL53L1X_chip_id[6]), 
         .Z(n37943)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i27267_3_lut.init = 16'hc8c8;
    PFUMX i167_adj_199 (.BLUT(n47989), .ALUT(n49085), .C0(tx_word_index[3]), 
          .Z(n117));
    PFUMX i40195 (.BLUT(n51042), .ALUT(n51041), .C0(\tx_byte_index[0] ), 
          .Z(n51043));
    L6MUX21 i169_adj_200 (.D0(n108_adj_5152), .D1(n117_adj_5153), .SD(n49682), 
            .Z(n123));
    L6MUX21 i169_adj_201 (.D0(n108_adj_5155), .D1(n117_adj_5156), .SD(n49682), 
            .Z(n123_adj_5157));
    L6MUX21 i25115 (.D0(n108_adj_5158), .D1(n117_adj_5159), .SD(n49682), 
            .Z(n37));
    LUT4 i39093_3_lut (.A(n2147[6]), .B(n37965), .C(\tx_byte_index[0] ), 
         .Z(n49483)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(96[17:30])
    defparam i39093_3_lut.init = 16'hcaca;
    PFUMX i167_adj_202 (.BLUT(n47990), .ALUT(n48928), .C0(tx_word_index[3]), 
          .Z(n117_adj_5159));
    LUT4 led_data_1__bdd_4_lut (.A(\led_data[1] ), .B(\led_data[3] ), .C(\led_data[0] ), 
         .D(\led_data[2] ), .Z(n51289)) /* synthesis lut_function=(A ((C)+!B)+!A !((C+!(D))+!B)) */ ;
    defparam led_data_1__bdd_4_lut.init = 16'ha6a2;
    PFUMX i167_adj_203 (.BLUT(n47988), .ALUT(n48972), .C0(tx_word_index[3]), 
          .Z(n117_adj_5153));
    PFUMX i167_adj_204 (.BLUT(n47987), .ALUT(n121), .C0(tx_word_index[3]), 
          .Z(n117_adj_5156));
    LUT4 i37622_3_lut (.A(state[3]), .B(\state[5] ), .C(state[8]), .Z(n15)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam i37622_3_lut.init = 16'h0101;
    LUT4 i37468_3_lut (.A(state[8]), .B(state[3]), .C(next_state_9__N_4541[6]), 
         .Z(n3_adj_5160)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam i37468_3_lut.init = 16'h0101;
    L6MUX21 i25128 (.D0(n108_adj_5161), .D1(n117_adj_5162), .SD(n49682), 
            .Z(n39_adj_5147));
    LUT4 i39223_3_lut (.A(n3_adj_5160), .B(n15), .C(state[4]), .Z(n17)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(218[13] 230[20])
    defparam i39223_3_lut.init = 16'hcaca;
    PFUMX i41036 (.BLUT(n51351), .ALUT(n52715), .C0(\tx_word_index[1] ), 
          .Z(n52716));
    LUT4 VL53L1X_chip_id_5__bdd_3_lut_4_lut (.A(VL53L1X_chip_id[0]), .B(VL53L1X_chip_id[1]), 
         .C(VL53L1X_chip_id[2]), .D(VL53L1X_chip_id[3]), .Z(n51008)) /* synthesis lut_function=(A (B)+!A !(B (D)+!B !(C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(237[13] 255[20])
    defparam VL53L1X_chip_id_5__bdd_3_lut_4_lut.init = 16'h98cc;
    PFUMX i167_adj_205 (.BLUT(n47986), .ALUT(n121_adj_5163), .C0(tx_word_index[3]), 
          .Z(n117_adj_5162));
    LUT4 mux_268_Mux_0_i15_3_lut_4_lut (.A(VL53L1X_chip_id[4]), .B(VL53L1X_chip_id[6]), 
         .C(VL53L1X_chip_id[5]), .D(VL53L1X_chip_id[7]), .Z(n2019[0])) /* synthesis lut_function=(!(A (B (D)+!B (C (D)))+!A !(B (D)+!B (C (D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(237[13] 255[20])
    defparam mux_268_Mux_0_i15_3_lut_4_lut.init = 16'h56aa;
    LUT4 i4_4_lut (.A(state[8]), .B(next_state_9__N_4571[5]), .C(n52451), 
         .D(n49291), .Z(next_state_9__N_4478[9])) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i4_4_lut.init = 16'h0002;
    LUT4 z_linear_velocity_13__bdd_3_lut_4_lut (.A(\z_linear_velocity[8] ), 
         .B(\z_linear_velocity[9] ), .C(\z_linear_velocity[10] ), .D(\z_linear_velocity[11] ), 
         .Z(n51015)) /* synthesis lut_function=(A (B)+!A !(B (D)+!B !(C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(237[13] 255[20])
    defparam z_linear_velocity_13__bdd_3_lut_4_lut.init = 16'h98cc;
    PFUMX i164 (.BLUT(n47968), .ALUT(n27741), .C0(tx_word_index[2]), .Z(n108));
    LUT4 n1_bdd_4_lut (.A(n1_adj_5106), .B(\tx_byte_index[1] ), .C(n53527), 
         .D(tx_byte_index[2]), .Z(n53871)) /* synthesis lut_function=(A (B (C (D))+!B (C+!(D)))+!A (C (D))) */ ;
    defparam n1_bdd_4_lut.init = 16'hf022;
    L6MUX21 i168 (.D0(n25957), .D1(n48295), .SD(tx_word_index[2]), .Z(n48486));
    PFUMX i40186 (.BLUT(n51028), .ALUT(n51027), .C0(\tx_byte_index[0] ), 
          .Z(n51029));
    L6MUX21 i168_adj_206 (.D0(n38452), .D1(n38456), .SD(n52407), .Z(n38458));
    LUT4 i2_4_lut_adj_207 (.A(n52255), .B(n52179), .C(n41_adj_5149), .D(n27735), 
         .Z(n48731)) /* synthesis lut_function=(A ((D)+!B)+!A ((C+(D))+!B)) */ ;
    defparam i2_4_lut_adj_207.init = 16'hff73;
    PFUMX i40791 (.BLUT(n51974), .ALUT(n51972), .C0(\tx_byte_index[1] ), 
          .Z(n51975));
    LUT4 i3_4_lut_adj_208 (.A(tx_word_index[7]), .B(tx_word_index[5]), .C(tx_word_index[6]), 
         .D(tx_word_index[3]), .Z(n47335)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(237[13] 255[20])
    defparam i3_4_lut_adj_208.init = 16'hfffe;
    LUT4 i1_4_lut_adj_209 (.A(n52240), .B(n81), .C(n52383), .D(tx_byte_index[2]), 
         .Z(n27735)) /* synthesis lut_function=(A (B (C+!(D)))+!A (B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(226[60:96])
    defparam i1_4_lut_adj_209.init = 16'hc088;
    LUT4 i1_2_lut_adj_210 (.A(n7_adj_5164), .B(n47552), .Z(next_state_9__N_4478[8])) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(218[13] 230[20])
    defparam i1_2_lut_adj_210.init = 16'h4444;
    LUT4 i19_1_lut_rep_506 (.A(tx_byte_index[2]), .Z(n52442)) /* synthesis lut_function=(!(A)) */ ;
    defparam i19_1_lut_rep_506.init = 16'h5555;
    LUT4 n48679_bdd_4_lut (.A(n43271), .B(\tx_byte_index[1] ), .C(yaw_val[1]), 
         .D(yaw_val[2]), .Z(n51316)) /* synthesis lut_function=(A (B+(D))+!A (B+(C (D)))) */ ;
    defparam n48679_bdd_4_lut.init = 16'hfecc;
    LUT4 n43228_bdd_4_lut (.A(n52390), .B(\tx_byte_index[1] ), .C(\VL53L1X_range_mm[6] ), 
         .D(\VL53L1X_range_mm[5] ), .Z(n50806)) /* synthesis lut_function=(A (B+(D))+!A (B+!((D)+!C))) */ ;
    defparam n43228_bdd_4_lut.init = 16'heedc;
    LUT4 n51322_bdd_3_lut_3_lut (.A(tx_byte_index[2]), .B(n34534), .C(n51322), 
         .Z(n51323)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam n51322_bdd_3_lut_3_lut.init = 16'he4e4;
    LUT4 i3_4_lut_adj_211 (.A(\tx_byte_index[0] ), .B(\tx_byte_index[1] ), 
         .C(tx_byte_index[2]), .D(tx_byte_index[3]), .Z(n7_adj_5164)) /* synthesis lut_function=(A+(B+(C+!(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(226[60:96])
    defparam i3_4_lut_adj_211.init = 16'hfeff;
    LUT4 n48676_bdd_3_lut (.A(n48676), .B(n27_adj_5165), .C(\tx_byte_index[0] ), 
         .Z(n51319)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n48676_bdd_3_lut.init = 16'hcaca;
    LUT4 i6_4_lut (.A(n52453), .B(n12), .C(state[7]), .D(\state[6] ), 
         .Z(n47552)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;
    defparam i6_4_lut.init = 16'h0040;
    LUT4 i5_4_lut_adj_212 (.A(next_state_9__N_4551[6]), .B(n52451), .C(n36607), 
         .D(n52342), .Z(n12)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i5_4_lut_adj_212.init = 16'h0002;
    LUT4 i38690_3_lut_3_lut (.A(tx_byte_index[2]), .B(n18), .C(n49484), 
         .Z(n49485)) /* synthesis lut_function=(A (C)+!A (B)) */ ;
    defparam i38690_3_lut_3_lut.init = 16'he4e4;
    LUT4 i1_2_lut_adj_213 (.A(state[4]), .B(\state[5] ), .Z(n36607)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam i1_2_lut_adj_213.init = 16'heeee;
    PFUMX i15483 (.BLUT(n49376), .ALUT(n49377), .C0(n49697), .Z(n25957));
    PFUMX i40178 (.BLUT(n51016), .ALUT(n51015), .C0(\tx_byte_index[0] ), 
          .Z(n51017));
    LUT4 i26107_3_lut (.A(latched_pitch[1]), .B(latched_pitch[3]), .C(latched_pitch[2]), 
         .Z(n1524[6])) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(237[13] 255[20])
    defparam i26107_3_lut.init = 16'hc8c8;
    LUT4 n50855_bdd_4_lut (.A(n14_adj_5166), .B(\tx_byte_index[1] ), .C(yaw_val[5]), 
         .D(yaw_val[7]), .Z(n51321)) /* synthesis lut_function=(A (B+(C+(D)))+!A (B+!((D)+!C))) */ ;
    defparam n50855_bdd_4_lut.init = 16'heefc;
    PFUMX i164_adj_214 (.BLUT(n47967), .ALUT(n27743), .C0(tx_word_index[2]), 
          .Z(n108_adj_5150));
    PFUMX i164_adj_215 (.BLUT(n47969), .ALUT(n27742), .C0(tx_word_index[2]), 
          .Z(n108_adj_5158));
    PFUMX i166 (.BLUT(n5_adj_5140), .ALUT(n25955), .C0(\tx_word_index[1] ), 
          .Z(n48295));
    LUT4 i26566_2_lut_rep_498 (.A(tx_word_index[5]), .B(tx_word_index[6]), 
         .Z(n52434)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(237[13] 255[20])
    defparam i26566_2_lut_rep_498.init = 16'heeee;
    LUT4 n12_bdd_4_lut (.A(n12_adj_5167), .B(\tx_byte_index[0] ), .C(\tx_byte_index[1] ), 
         .D(n50824), .Z(n51324)) /* synthesis lut_function=(A (B+(C+(D)))+!A !(B+!(C+(D)))) */ ;
    defparam n12_bdd_4_lut.init = 16'hbbb8;
    LUT4 i1_2_lut_3_lut_4_lut_adj_216 (.A(tx_word_index[5]), .B(tx_word_index[6]), 
         .C(n123_adj_5157), .D(tx_word_index[7]), .Z(n27651)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(237[13] 255[20])
    defparam i1_2_lut_3_lut_4_lut_adj_216.init = 16'h0010;
    LUT4 i86_2_lut_rep_319_3_lut (.A(tx_word_index[5]), .B(tx_word_index[6]), 
         .C(tx_word_index[7]), .Z(n52255)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(237[13] 255[20])
    defparam i86_2_lut_rep_319_3_lut.init = 16'hfefe;
    LUT4 i3_4_lut_adj_217 (.A(state[4]), .B(n22_adj_5168), .C(n38171), 
         .D(state[7]), .Z(next_state_9__N_4478[6])) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i3_4_lut_adj_217.init = 16'h0004;
    LUT4 n34657_bdd_4_lut_40712_4_lut_rep_443_3_lut (.A(\tx_word_index[1] ), 
         .B(tx_word_index[0]), .C(tx_word_index[2]), .Z(n52379)) /* synthesis lut_function=(A+!(B+(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(371[42:62])
    defparam n34657_bdd_4_lut_40712_4_lut_rep_443_3_lut.init = 16'habab;
    LUT4 i166_4_lut_4_lut_4_lut (.A(tx_word_index[2]), .B(n25927), .C(n38373), 
         .D(n52398), .Z(n114)) /* synthesis lut_function=(!(A ((D)+!C)+!A ((D)+!B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(371[42:62])
    defparam i166_4_lut_4_lut_4_lut.init = 16'h00e4;
    LUT4 i33_4_lut (.A(next_state_9__N_4541[6]), .B(\state[6] ), .C(\state[5] ), 
         .D(next_state_9__N_4551[6]), .Z(n22_adj_5168)) /* synthesis lut_function=(!(A (B (C+!(D))+!B !(C))+!A ((C+!(D))+!B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(218[13] 230[20])
    defparam i33_4_lut.init = 16'h2c20;
    LUT4 i4_4_lut_adj_218 (.A(n52257), .B(state[7]), .C(\state[6] ), .D(n6_adj_5169), 
         .Z(next_state_9__N_4478[5])) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i4_4_lut_adj_218.init = 16'h0100;
    LUT4 i27280_3_lut (.A(latched_pitch[5]), .B(latched_pitch[7]), .C(latched_pitch[6]), 
         .Z(n37957)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i27280_3_lut.init = 16'hc8c8;
    PFUMX i166_adj_219 (.BLUT(n38444), .ALUT(n38454), .C0(n52378), .Z(n38456));
    LUT4 i1_2_lut_adj_220 (.A(n7_adj_5164), .B(n47552), .Z(next_state_9__N_4478[4])) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(218[13] 230[20])
    defparam i1_2_lut_adj_220.init = 16'h8888;
    LUT4 i1_2_lut_3_lut_adj_221 (.A(\VL53L1X_range_mm[9] ), .B(\VL53L1X_range_mm[10] ), 
         .C(\VL53L1X_range_mm[11] ), .Z(n5)) /* synthesis lut_function=(A (C)+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(155[9:25])
    defparam i1_2_lut_3_lut_adj_221.init = 16'he0e0;
    PFUMX i164_adj_222 (.BLUT(n47965), .ALUT(n91), .C0(tx_word_index[2]), 
          .Z(n108_adj_5155));
    LUT4 n53077_bdd_3_lut_41267 (.A(n53077), .B(n53076), .C(tx_word_index[2]), 
         .Z(n53078)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n53077_bdd_3_lut_41267.init = 16'hcaca;
    LUT4 i1_2_lut_adj_223 (.A(\state[2] ), .B(n45947), .Z(n6_adj_5169)) /* synthesis lut_function=(!(A+!(B))) */ ;
    defparam i1_2_lut_adj_223.init = 16'h4444;
    LUT4 i2_4_lut_adj_224 (.A(\state[5] ), .B(n4_adj_5170), .C(\state[6] ), 
         .D(n27995), .Z(n47346)) /* synthesis lut_function=(A (B)+!A (B+!((D)+!C))) */ ;
    defparam i2_4_lut_adj_224.init = 16'hccdc;
    LUT4 i1_4_lut_adj_225 (.A(n37479), .B(state[7]), .C(n52453), .D(n52206), 
         .Z(n4_adj_5170)) /* synthesis lut_function=(!(A ((C+(D))+!B))) */ ;
    defparam i1_4_lut_adj_225.init = 16'h555d;
    LUT4 i15490_4_lut_4_lut (.A(tx_byte_index[2]), .B(n52383), .C(n52240), 
         .D(n34504), .Z(n25964)) /* synthesis lut_function=(A (B+(D))+!A (C)) */ ;
    defparam i15490_4_lut_4_lut.init = 16'hfad8;
    LUT4 i1_2_lut_rep_304_2_lut (.A(\tx_byte_index[1] ), .B(n1_adj_5106), 
         .Z(n52240)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam i1_2_lut_rep_304_2_lut.init = 16'h4444;
    LUT4 i1_4_lut_adj_226 (.A(\tx_byte_index[1] ), .B(VL53L1X_firm_rdy[0]), 
         .C(VL53L1X_firm_rdy[2]), .D(n48161), .Z(n27_adj_5122)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(265[13] 275[20])
    defparam i1_4_lut_adj_226.init = 16'hfaea;
    LUT4 i2_4_lut_4_lut (.A(\tx_byte_index[1] ), .B(n41683), .C(\amc_debug[6] ), 
         .D(\amc_debug[5] ), .Z(n48537)) /* synthesis lut_function=(!(A+!(B (C)+!B (C (D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam i2_4_lut_4_lut.init = 16'h5040;
    LUT4 n51202_bdd_4_lut_4_lut (.A(\tx_byte_index[1] ), .B(\tx_word_index[1] ), 
         .C(n51201), .D(n51202), .Z(n52166)) /* synthesis lut_function=(A+!(B (C)+!B (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam n51202_bdd_4_lut_4_lut.init = 16'haebf;
    LUT4 i3_3_lut_4_lut_4_lut_4_lut (.A(\tx_byte_index[1] ), .B(n18), .C(n81), 
         .D(tx_byte_index[2]), .Z(n49126)) /* synthesis lut_function=(!(A+(((D)+!C)+!B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam i3_3_lut_4_lut_4_lut_4_lut.init = 16'h0040;
    LUT4 n28_bdd_4_lut_4_lut (.A(\tx_byte_index[1] ), .B(n50977), .C(n51159), 
         .D(\tx_word_index[1] ), .Z(n51353)) /* synthesis lut_function=(!(A+!(B (C+(D))+!B !((D)+!C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam n28_bdd_4_lut_4_lut.init = 16'h4450;
    LUT4 i2_4_lut_4_lut_adj_227 (.A(\tx_byte_index[1] ), .B(n34474), .C(VL53L1X_data_rdy[5]), 
         .D(VL53L1X_data_rdy[6]), .Z(n48742)) /* synthesis lut_function=(!(A+!(B (D)+!B (C (D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam i2_4_lut_4_lut_adj_227.init = 16'h5400;
    LUT4 i2_4_lut_4_lut_adj_228 (.A(\tx_byte_index[1] ), .B(n52328), .C(latched_pitch[6]), 
         .D(latched_pitch[4]), .Z(n48692)) /* synthesis lut_function=(!(A+!(B (C)+!B (C (D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam i2_4_lut_4_lut_adj_228.init = 16'h5040;
    LUT4 i26137_2_lut_2_lut (.A(\tx_byte_index[1] ), .B(n1), .Z(n20)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam i26137_2_lut_2_lut.init = 16'h4444;
    LUT4 i43_4_lut_3_lut (.A(\tx_byte_index[1] ), .B(n51289), .C(\tx_byte_index[0] ), 
         .Z(n23)) /* synthesis lut_function=(!(A (C)+!A !(B (C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam i43_4_lut_3_lut.init = 16'h4a4a;
    LUT4 n51581_bdd_4_lut_4_lut (.A(\tx_byte_index[1] ), .B(\tx_byte_index[0] ), 
         .C(n51580), .D(n51581), .Z(n34534)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam n51581_bdd_4_lut_4_lut.init = 16'h5140;
    LUT4 i25986_2_lut_2_lut (.A(\tx_byte_index[1] ), .B(n37975), .Z(n6_adj_5141)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam i25986_2_lut_2_lut.init = 16'h4444;
    LUT4 i1_2_lut_2_lut (.A(\tx_byte_index[1] ), .B(\i2c_device_driver_return_state[4] ), 
         .Z(n13)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam i1_2_lut_2_lut.init = 16'h4444;
    LUT4 i38681_3_lut_4_lut_4_lut_4_lut (.A(\tx_byte_index[1] ), .B(n1_adj_5106), 
         .C(n50721), .D(tx_byte_index[2]), .Z(n49476)) /* synthesis lut_function=(A (C (D))+!A (B (C+!(D))+!B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam i38681_3_lut_4_lut_4_lut_4_lut.init = 16'hf044;
    LUT4 n11_bdd_4_lut_4_lut (.A(\tx_byte_index[1] ), .B(tx_word_index[0]), 
         .C(n19), .D(n51273), .Z(n52158)) /* synthesis lut_function=(A (B (C))+!A (B (C)+!B (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam n11_bdd_4_lut_4_lut.init = 16'hd1c0;
    LUT4 i1_4_lut_4_lut_adj_229 (.A(\tx_byte_index[1] ), .B(n52419), .C(VL53L1X_data_rdy[7]), 
         .D(VL53L1X_data_rdy[4]), .Z(n39)) /* synthesis lut_function=(!(A+(B (C (D)+!C !(D))+!B !(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam i1_4_lut_4_lut_adj_229.init = 16'h1540;
    PFUMX i164_adj_230 (.BLUT(n47966), .ALUT(n27740), .C0(tx_word_index[2]), 
          .Z(n108_adj_5152));
    LUT4 i2_4_lut_4_lut_adj_231 (.A(\tx_byte_index[1] ), .B(n52422), .C(yaw_val[6]), 
         .D(yaw_val[4]), .Z(n48679)) /* synthesis lut_function=(!(A+!(B (C)+!B (C (D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam i2_4_lut_4_lut_adj_231.init = 16'h5040;
    LUT4 gnd_bdd_2_lut_40015_2_lut (.A(\tx_byte_index[1] ), .B(n50719), 
         .Z(n50720)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam gnd_bdd_2_lut_40015_2_lut.init = 16'h4444;
    LUT4 n43228_bdd_4_lut_40041_4_lut (.A(\tx_byte_index[1] ), .B(\VL53L1X_range_mm[1] ), 
         .C(\VL53L1X_range_mm[2] ), .D(n52388), .Z(n50805)) /* synthesis lut_function=(!(A+!(B (D)+!B !((D)+!C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam n43228_bdd_4_lut_40041_4_lut.init = 16'h4410;
    LUT4 i2_4_lut_then_4_lut (.A(\state[5] ), .B(state[9]), .C(state[3]), 
         .D(next_state_9__N_4541[6]), .Z(n52511)) /* synthesis lut_function=(!(A+(B+(C+!(D))))) */ ;
    defparam i2_4_lut_then_4_lut.init = 16'h0100;
    LUT4 n34481_bdd_4_lut_40074_4_lut (.A(\tx_byte_index[1] ), .B(VL53L1X_data_rdy[2]), 
         .C(VL53L1X_data_rdy[1]), .D(n52389), .Z(n50858)) /* synthesis lut_function=(!(A+!(B (C (D)+!C !(D))+!B (C (D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam n34481_bdd_4_lut_40074_4_lut.init = 16'h5004;
    PFUMX i164_adj_232 (.BLUT(n48823), .ALUT(n48839), .C0(tx_word_index[2]), 
          .Z(n108_adj_5161));
    LUT4 i38631_4_lut_4_lut (.A(\tx_byte_index[1] ), .B(tx_byte_index[2]), 
         .C(n43217), .D(n38325), .Z(n49426)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam i38631_4_lut_4_lut.init = 16'h7340;
    LUT4 i38632_4_lut_4_lut (.A(\tx_byte_index[1] ), .B(tx_byte_index[2]), 
         .C(n43303), .D(n38329), .Z(n49427)) /* synthesis lut_function=(!(A (B+!(D))+!A !(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam i38632_4_lut_4_lut.init = 16'h7340;
    LUT4 i2_4_lut_4_lut_adj_233 (.A(\tx_byte_index[1] ), .B(n48147), .C(VL53L1X_firm_rdy[6]), 
         .D(VL53L1X_firm_rdy[4]), .Z(n48706)) /* synthesis lut_function=(!(A+!(B (C)+!B (C (D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam i2_4_lut_4_lut_adj_233.init = 16'h5040;
    LUT4 i1_4_lut_4_lut_adj_234 (.A(\tx_byte_index[1] ), .B(latched_pitch[7]), 
         .C(n14_adj_5145), .D(latched_pitch[4]), .Z(n13_adj_5127)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam i1_4_lut_4_lut_adj_234.init = 16'h5140;
    LUT4 n28_bdd_3_lut (.A(n28), .B(n12_adj_5171), .C(\tx_byte_index[0] ), 
         .Z(n51351)) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;
    defparam n28_bdd_3_lut.init = 16'hcaca;
    LUT4 i2_3_lut_3_lut (.A(\tx_byte_index[1] ), .B(n47964), .C(n99_adj_5125), 
         .Z(n48823)) /* synthesis lut_function=(!(A+!(B (C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam i2_3_lut_3_lut.init = 16'h4040;
    LUT4 gnd_bdd_2_lut_40551_2_lut (.A(\tx_byte_index[1] ), .B(n51610), 
         .Z(n51611)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam gnd_bdd_2_lut_40551_2_lut.init = 16'h4444;
    LUT4 n26269_bdd_4_lut_4_lut (.A(tx_word_index[2]), .B(n49482), .C(\tx_byte_index[1] ), 
         .D(n26269), .Z(n51627)) /* synthesis lut_function=(A (B+(C))+!A (C+(D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(371[42:62])
    defparam n26269_bdd_4_lut_4_lut.init = 16'hfdf8;
    LUT4 i1_4_lut_4_lut_adj_235 (.A(\tx_byte_index[1] ), .B(swa_swb_val[7]), 
         .C(n14_adj_5146), .D(swa_swb_val[4]), .Z(n13_adj_5128)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam i1_4_lut_4_lut_adj_235.init = 16'h5140;
    LUT4 gnd_bdd_2_lut_40650_2_lut (.A(\tx_byte_index[1] ), .B(n51747), 
         .Z(n51748)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam gnd_bdd_2_lut_40650_2_lut.init = 16'h4444;
    LUT4 i1_4_lut_adj_236 (.A(\tx_byte_index[1] ), .B(\amc_debug[1] ), .C(\amc_debug[2] ), 
         .D(n41688), .Z(n71)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam i1_4_lut_adj_236.init = 16'hfaea;
    LUT4 i1_4_lut_4_lut_4_lut_adj_237 (.A(\tx_byte_index[1] ), .B(throttle_val[1]), 
         .C(n52429), .D(throttle_val[2]), .Z(n12_adj_5167)) /* synthesis lut_function=(!(A+!(B (C)+!B !(C+!(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam i1_4_lut_4_lut_4_lut_adj_237.init = 16'h4140;
    LUT4 n43271_bdd_4_lut_40071_4_lut (.A(\tx_byte_index[1] ), .B(yaw_val[1]), 
         .C(yaw_val[2]), .D(n43271), .Z(n50855)) /* synthesis lut_function=(!(A+!(B (D)+!B !((D)+!C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam n43271_bdd_4_lut_40071_4_lut.init = 16'h4410;
    LUT4 gnd_bdd_2_lut_40643_2_lut (.A(\tx_byte_index[1] ), .B(n51743), 
         .Z(n51744)) /* synthesis lut_function=(!(A+!(B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam gnd_bdd_2_lut_40643_2_lut.init = 16'h4444;
    L6MUX21 i38917 (.D0(n49710), .D1(n49711), .SD(tx_word_index[0]), .Z(n49712));
    LUT4 i2_4_lut_4_lut_adj_238 (.A(\tx_byte_index[1] ), .B(n52437), .C(throttle_val[6]), 
         .D(throttle_val[4]), .Z(n48676)) /* synthesis lut_function=(!(A+!(B (C)+!B (C (D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam i2_4_lut_4_lut_adj_238.init = 16'h5040;
    LUT4 i1_4_lut_4_lut_adj_239 (.A(\tx_byte_index[1] ), .B(latched_pitch[3]), 
         .C(n36752), .D(latched_pitch[1]), .Z(n12_adj_5171)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam i1_4_lut_4_lut_adj_239.init = 16'h5140;
    LUT4 i1_4_lut_4_lut_adj_240 (.A(\tx_byte_index[1] ), .B(\latched_roll[7] ), 
         .C(n14_adj_5144), .D(\latched_roll[4] ), .Z(n13_adj_5126)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam i1_4_lut_4_lut_adj_240.init = 16'h5140;
    LUT4 n41683_bdd_4_lut_40364_4_lut (.A(\tx_byte_index[1] ), .B(\amc_debug[1] ), 
         .C(\amc_debug[2] ), .D(n41688), .Z(n51326)) /* synthesis lut_function=(!(A+!(B (D)+!B !((D)+!C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam n41683_bdd_4_lut_40364_4_lut.init = 16'h4410;
    LUT4 i2_3_lut_3_lut_rep_507 (.A(\tx_byte_index[1] ), .B(tx_byte_index[3]), 
         .C(tx_byte_index[2]), .Z(n52443)) /* synthesis lut_function=((B+(C))+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam i2_3_lut_3_lut_rep_507.init = 16'hfdfd;
    LUT4 i2_4_lut_else_4_lut (.A(\state[5] ), .B(next_state_9__N_4531[5]), 
         .C(state[9]), .D(state[3]), .Z(n52510)) /* synthesis lut_function=(!(A+(B ((D)+!C)+!B (C (D)+!C !(D))))) */ ;
    defparam i2_4_lut_else_4_lut.init = 16'h0150;
    LUT4 i27709_3_lut_4_lut_4_lut (.A(\tx_byte_index[1] ), .B(tx_byte_index[3]), 
         .C(tx_byte_index[2]), .D(n38373), .Z(n38444)) /* synthesis lut_function=(A (B+(C))+!A (B+(D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam i27709_3_lut_4_lut_4_lut.init = 16'hfdec;
    LUT4 i27716_3_lut_4_lut_4_lut (.A(\tx_byte_index[1] ), .B(tx_byte_index[3]), 
         .C(tx_byte_index[2]), .D(n25927), .Z(n38454)) /* synthesis lut_function=(A (B+(C))+!A (B+(D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam i27716_3_lut_4_lut_4_lut.init = 16'hfdec;
    LUT4 i27697_3_lut_4_lut_4_lut (.A(\tx_byte_index[1] ), .B(tx_byte_index[3]), 
         .C(tx_byte_index[2]), .D(n24), .Z(n38432)) /* synthesis lut_function=(A (B+(C))+!A (B+(D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam i27697_3_lut_4_lut_4_lut.init = 16'hfdec;
    LUT4 mux_204_Mux_1_i14_4_lut_3_lut (.A(latched_pitch[4]), .B(latched_pitch[5]), 
         .C(latched_pitch[6]), .Z(n14_adj_5172)) /* synthesis lut_function=(A (B)+!A !(B+!(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(237[13] 255[20])
    defparam mux_204_Mux_1_i14_4_lut_3_lut.init = 16'h9898;
    LUT4 i15458_4_lut_4_lut (.A(\tx_word_index[1] ), .B(tx_byte_index[2]), 
         .C(n50886), .D(n49435), .Z(n25927)) /* synthesis lut_function=(A (C)+!A (B (D)+!B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(371[42:62])
    defparam i15458_4_lut_4_lut.init = 16'hf4b0;
    PFUMX i41510 (.BLUT(n53558), .ALUT(n53557), .C0(\tx_byte_index[0] ), 
          .Z(n53559));
    L6MUX21 i38606 (.D0(n49399), .D1(n49400), .SD(tx_word_index[0]), .Z(n49401));
    L6MUX21 i41492 (.D0(n53871), .D1(n53526), .SD(tx_word_index[0]), .Z(n49448));
    PFUMX i41488 (.BLUT(n53525), .ALUT(n53524), .C0(\tx_byte_index[0] ), 
          .Z(n53526));
    LUT4 i1_4_lut_adj_241 (.A(\tx_byte_index[1] ), .B(latched_pitch[5]), 
         .C(n14_adj_5172), .D(latched_pitch[7]), .Z(n28)) /* synthesis lut_function=(A+(B (C+!(D))+!B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(265[13] 275[20])
    defparam i1_4_lut_adj_241.init = 16'hfaee;
    PFUMX i39984 (.BLUT(n50675), .ALUT(n50674), .C0(\tx_byte_index[0] ), 
          .Z(n50676));
    PFUMX i161 (.BLUT(n38432), .ALUT(n38447), .C0(tx_word_index[0]), .Z(n38452));
    L6MUX21 i41413 (.D0(n53397), .D1(n53395), .SD(tx_word_index[0]), .Z(n53398));
    PFUMX i41411 (.BLUT(n53396), .ALUT(n51135), .C0(\tx_byte_index[0] ), 
          .Z(n53397));
    PFUMX i41409 (.BLUT(n53394), .ALUT(n52541), .C0(\tx_byte_index[0] ), 
          .Z(n53395));
    PFUMX i40644 (.BLUT(n51748), .ALUT(n51746), .C0(\tx_byte_index[0] ), 
          .Z(n51749));
    L6MUX21 i41404 (.D0(n53384), .D1(n53382), .SD(tx_word_index[0]), .Z(n53385));
    PFUMX i41400 (.BLUT(n53381), .ALUT(n50715), .C0(\tx_byte_index[0] ), 
          .Z(n53382));
    PFUMX i41402 (.BLUT(n53383), .ALUT(n25), .C0(\tx_byte_index[0] ), 
          .Z(n53384));
    PFUMX i35 (.BLUT(n20_adj_5148), .ALUT(n17), .C0(n36607), .Z(n45947));
    PFUMX i40640 (.BLUT(n51744), .ALUT(n51742), .C0(\tx_byte_index[0] ), 
          .Z(n51745));
    PFUMX i38915 (.BLUT(n49706), .ALUT(n52167), .C0(tx_byte_index[2]), 
          .Z(n49710));
    PFUMX i38916 (.BLUT(n49708), .ALUT(n49709), .C0(tx_byte_index[2]), 
          .Z(n49711));
    L6MUX21 i38945 (.D0(n49738), .D1(n49739), .SD(\tx_word_index[1] ), 
            .Z(n49740));
    LUT4 i1_2_lut_rep_258_3_lut_4_lut (.A(n52454), .B(n52294), .C(state[7]), 
         .D(n48129), .Z(n52194)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(366[17:29])
    defparam i1_2_lut_rep_258_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_4_lut_adj_242 (.A(n52194), .B(state[8]), .C(state[9]), 
         .D(n7), .Z(n64)) /* synthesis lut_function=(A (D)+!A (B ((D)+!C)+!B (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(366[17:29])
    defparam i1_2_lut_4_lut_adj_242.init = 16'hff04;
    LUT4 i39855_2_lut_3_lut (.A(n52180), .B(n52179), .C(n52196), .Z(next_adr_i_7__N_4470[0])) /* synthesis lut_function=(A+!(B (C))) */ ;
    defparam i39855_2_lut_3_lut.init = 16'hbfbf;
    LUT4 i1_2_lut_rep_259_3_lut_4_lut (.A(n48129), .B(n52295), .C(state[4]), 
         .D(n52454), .Z(n52195)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(299[17:22])
    defparam i1_2_lut_rep_259_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_515 (.A(state[3]), .B(\state[2] ), .Z(n52451)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam i1_2_lut_rep_515.init = 16'heeee;
    LUT4 i27371_3_lut (.A(yaw_val[5]), .B(yaw_val[7]), .C(yaw_val[6]), 
         .Z(n38059)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i27371_3_lut.init = 16'hc8c8;
    LUT4 i4888_1_lut (.A(\led_data[1] ), .Z(\led_data_out_7__N_1[2] )) /* synthesis lut_function=(!(A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(237[13] 255[20])
    defparam i4888_1_lut.init = 16'h5555;
    LUT4 i1_2_lut_rep_358_3_lut (.A(state[3]), .B(\state[2] ), .C(state[4]), 
         .Z(n52294)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam i1_2_lut_rep_358_3_lut.init = 16'hfefe;
    LUT4 i39815_2_lut_4_lut (.A(n52194), .B(state[8]), .C(state[9]), .D(n7), 
         .Z(sys_clk_enable_217)) /* synthesis lut_function=(!(A (D)+!A (B (C (D))+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(366[17:29])
    defparam i39815_2_lut_4_lut.init = 16'h04ff;
    LUT4 i1_2_lut_rep_308_3_lut_4_lut (.A(state[3]), .B(\state[2] ), .C(n52454), 
         .D(state[4]), .Z(n52244)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam i1_2_lut_rep_308_3_lut_4_lut.init = 16'hfffe;
    PFUMX i41324 (.BLUT(n34534), .ALUT(n53238), .C0(tx_byte_index[2]), 
          .Z(n53239));
    L6MUX21 i41322 (.D0(n53236), .D1(n53234), .SD(\tx_word_index[1] ), 
            .Z(n53237));
    LUT4 i1_2_lut_4_lut_adj_243 (.A(n52194), .B(state[8]), .C(state[9]), 
         .D(n7), .Z(n40212)) /* synthesis lut_function=(!(A (D)+!A (B ((D)+!C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(366[17:29])
    defparam i1_2_lut_4_lut_adj_243.init = 16'h00fb;
    PFUMX i41320 (.BLUT(n53235), .ALUT(n9499[1]), .C0(tx_word_index[0]), 
          .Z(n53236));
    LUT4 i1_2_lut_4_lut_adj_244 (.A(n52195), .B(state[3]), .C(\state[2] ), 
         .D(n15182), .Z(n48081)) /* synthesis lut_function=(A (D)+!A (B (D)+!B !(C+!(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam i1_2_lut_4_lut_adj_244.init = 16'hef00;
    LUT4 i27288_3_lut (.A(VL53L1X_firm_rdy[1]), .B(VL53L1X_firm_rdy[3]), 
         .C(VL53L1X_firm_rdy[2]), .Z(n37965)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i27288_3_lut.init = 16'hc8c8;
    PFUMX i41318 (.BLUT(n34534), .ALUT(n53233), .C0(tx_byte_index[2]), 
          .Z(n53234));
    LUT4 tx_byte_index_1__bdd_4_lut_40155 (.A(throttle_val[5]), .B(throttle_val[7]), 
         .C(throttle_val[4]), .D(throttle_val[6]), .Z(n50824)) /* synthesis lut_function=(A ((C)+!B)+!A !((C+!(D))+!B)) */ ;
    defparam tx_byte_index_1__bdd_4_lut_40155.init = 16'ha6a2;
    LUT4 i25643_3_lut (.A(VL53L1X_firm_rdy[5]), .B(VL53L1X_firm_rdy[7]), 
         .C(VL53L1X_firm_rdy[6]), .Z(n2147[6])) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(237[13] 255[20])
    defparam i25643_3_lut.init = 16'hc8c8;
    LUT4 i1_2_lut_rep_517 (.A(state[8]), .B(state[9]), .Z(n52453)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam i1_2_lut_rep_517.init = 16'heeee;
    LUT4 i37453_3_lut_4_lut (.A(n48129), .B(n52295), .C(state[0]), .D(state[1]), 
         .Z(n48229)) /* synthesis lut_function=(A+(B+(C (D)+!C !(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(299[17:22])
    defparam i37453_3_lut_4_lut.init = 16'hfeef;
    LUT4 i1_2_lut_rep_309_3_lut_4_lut (.A(state[8]), .B(state[9]), .C(n48129), 
         .D(state[7]), .Z(n52245)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam i1_2_lut_rep_309_3_lut_4_lut.init = 16'hfffe;
    LUT4 i1_4_lut_adj_245 (.A(\tx_byte_index[1] ), .B(throttle_val[1]), 
         .C(throttle_val[2]), .D(n52429), .Z(n27_adj_5165)) /* synthesis lut_function=(A+(B (C)+!B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam i1_4_lut_adj_245.init = 16'hfaea;
    LUT4 i27391_3_lut (.A(throttle_val[5]), .B(throttle_val[7]), .C(throttle_val[6]), 
         .Z(n38081)) /* synthesis lut_function=(A (B)+!A (B (C))) */ ;
    defparam i27391_3_lut.init = 16'hc8c8;
    LUT4 i1_2_lut_rep_359_3_lut (.A(state[8]), .B(state[9]), .C(state[7]), 
         .Z(n52295)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam i1_2_lut_rep_359_3_lut.init = 16'hfefe;
    LUT4 i1_2_lut_3_lut_adj_246 (.A(state[8]), .B(state[9]), .C(state[3]), 
         .Z(n37731)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam i1_2_lut_3_lut_adj_246.init = 16'hfefe;
    LUT4 state_9__I_0_i11_2_lut_rep_518 (.A(state[0]), .B(state[1]), .Z(n52454)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(373[17:24])
    defparam state_9__I_0_i11_2_lut_rep_518.init = 16'heeee;
    LUT4 i38489_2_lut_3_lut (.A(state[0]), .B(state[1]), .C(\state[2] ), 
         .Z(n49281)) /* synthesis lut_function=(A+(B+(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(373[17:24])
    defparam i38489_2_lut_3_lut.init = 16'hfefe;
    LUT4 mux_172_Mux_1_i14_4_lut_3_lut (.A(yaw_val[4]), .B(yaw_val[5]), 
         .C(yaw_val[6]), .Z(n14_adj_5166)) /* synthesis lut_function=(A (B)+!A !(B+!(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(237[13] 255[20])
    defparam mux_172_Mux_1_i14_4_lut_3_lut.init = 16'h9898;
    PFUMX i40104 (.BLUT(n50895), .ALUT(n18), .C0(n52442), .Z(n50896));
    LUT4 i1_2_lut_4_lut_4_lut (.A(tx_word_index[4]), .B(n52407), .C(n114), 
         .D(n99), .Z(n121_adj_5163)) /* synthesis lut_function=(!(A+!(B (C)+!B (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(227[46:89])
    defparam i1_2_lut_4_lut_4_lut.init = 16'h5140;
    PFUMX i40992 (.BLUT(n52597), .ALUT(n52598), .C0(\tx_byte_index[0] ), 
          .Z(n52599));
    LUT4 i4_4_lut_4_lut (.A(tx_word_index[4]), .B(n6_adj_5174), .C(tx_word_index[0]), 
         .D(n47335), .Z(next_state_9__N_4571[5])) /* synthesis lut_function=((B+((D)+!C))+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(227[46:89])
    defparam i4_4_lut_4_lut.init = 16'hffdf;
    PFUMX i40990 (.BLUT(n52594), .ALUT(n52595), .C0(\tx_byte_index[0] ), 
          .Z(n52596));
    L6MUX21 i40096 (.D0(n52160), .D1(n50882), .SD(n52375), .Z(n50886));
    PFUMX i40984 (.BLUT(n52585), .ALUT(n52586), .C0(\tx_byte_index[0] ), 
          .Z(n52587));
    PFUMX i40092 (.BLUT(n50881), .ALUT(n18), .C0(n52442), .Z(n50882));
    PFUMX i40972 (.BLUT(n52567), .ALUT(n52568), .C0(\tx_byte_index[0] ), 
          .Z(n34729));
    L6MUX21 i40562 (.D0(n51630), .D1(n51628), .SD(n52407), .Z(n51631));
    PFUMX i40558 (.BLUT(n34729), .ALUT(n51627), .C0(tx_byte_index[2]), 
          .Z(n51628));
    PFUMX i40560 (.BLUT(n51629), .ALUT(n9499[3]), .C0(tx_word_index[0]), 
          .Z(n51630));
    PFUMX i40968 (.BLUT(n52561), .ALUT(n52562), .C0(\tx_byte_index[0] ), 
          .Z(n52563));
    PFUMX i38605 (.BLUT(n3_adj_5111), .ALUT(n52168), .C0(tx_byte_index[2]), 
          .Z(n49400));
    PFUMX i40547 (.BLUT(n51613), .ALUT(n51611), .C0(\tx_byte_index[0] ), 
          .Z(n49411));
    PFUMX i38604 (.BLUT(n3_adj_5109), .ALUT(n52169), .C0(tx_byte_index[2]), 
          .Z(n49399));
    LUT4 i39732_2_lut_rep_439 (.A(tx_byte_index[2]), .B(tx_word_index[0]), 
         .Z(n52375)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(333[21] 354[28])
    defparam i39732_2_lut_rep_439.init = 16'hdddd;
    LUT4 i1_2_lut_2_lut_adj_247 (.A(\tx_word_index[1] ), .B(tx_word_index[2]), 
         .Z(n6_adj_5174)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(371[42:62])
    defparam i1_2_lut_2_lut_adj_247.init = 16'hdddd;
    LUT4 i39346_3_lut_4_lut (.A(tx_byte_index[2]), .B(tx_word_index[0]), 
         .C(n49476), .D(n51745), .Z(n25959)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(333[21] 354[28])
    defparam i39346_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i40948 (.BLUT(n52531), .ALUT(n52532), .C0(\tx_word_index[1] ), 
          .Z(n81));
    LUT4 i39310_3_lut_4_lut (.A(tx_byte_index[2]), .B(tx_word_index[0]), 
         .C(n25964), .D(n51749), .Z(n25965)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(333[21] 354[28])
    defparam i39310_3_lut_4_lut.init = 16'hf2d0;
    PFUMX i40946 (.BLUT(n52528), .ALUT(n52529), .C0(\tx_byte_index[0] ), 
          .Z(n52530));
    LUT4 i1_4_lut_adj_248 (.A(\tx_byte_index[1] ), .B(\i2c_device_driver_return_state[0] ), 
         .C(\i2c_device_driver_return_state[3] ), .D(n52457), .Z(n27_adj_5107)) /* synthesis lut_function=(A+!(B (C (D))+!B !(C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam i1_4_lut_adj_248.init = 16'hbeee;
    LUT4 n50897_bdd_3_lut_4_lut (.A(tx_byte_index[2]), .B(tx_word_index[0]), 
         .C(n50896), .D(n50897), .Z(n25919)) /* synthesis lut_function=(A (B (C)+!B (D))+!A (C)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(333[21] 354[28])
    defparam n50897_bdd_3_lut_4_lut.init = 16'hf2d0;
    FD1P3IX tx_word_index_6624__i7 (.D(n8[7]), .SP(sys_clk_enable_217), 
            .CD(n40212), .CK(sys_clk), .Q(tx_word_index[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(371[42:62])
    defparam tx_word_index_6624__i7.GSR = "ENABLED";
    FD1P3IX tx_word_index_6624__i6 (.D(n8[6]), .SP(sys_clk_enable_217), 
            .CD(n40212), .CK(sys_clk), .Q(tx_word_index[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(371[42:62])
    defparam tx_word_index_6624__i6.GSR = "ENABLED";
    FD1P3IX tx_word_index_6624__i5 (.D(n8[5]), .SP(sys_clk_enable_217), 
            .CD(n40212), .CK(sys_clk), .Q(tx_word_index[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(371[42:62])
    defparam tx_word_index_6624__i5.GSR = "ENABLED";
    FD1P3IX tx_word_index_6624__i4 (.D(n8[4]), .SP(sys_clk_enable_217), 
            .CD(n40212), .CK(sys_clk), .Q(tx_word_index[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(371[42:62])
    defparam tx_word_index_6624__i4.GSR = "ENABLED";
    FD1P3IX tx_word_index_6624__i3 (.D(n8[3]), .SP(sys_clk_enable_217), 
            .CD(n40212), .CK(sys_clk), .Q(tx_word_index[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(371[42:62])
    defparam tx_word_index_6624__i3.GSR = "ENABLED";
    FD1P3IX tx_word_index_6624__i2 (.D(n8[2]), .SP(sys_clk_enable_217), 
            .CD(n40212), .CK(sys_clk), .Q(tx_word_index[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(371[42:62])
    defparam tx_word_index_6624__i2.GSR = "ENABLED";
    FD1P3IX tx_word_index_6624__i1 (.D(n8[1]), .SP(sys_clk_enable_217), 
            .CD(n40212), .CK(sys_clk), .Q(\tx_word_index[1] )) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(371[42:62])
    defparam tx_word_index_6624__i1.GSR = "ENABLED";
    FD1P3IX tx_byte_index_6622__i3 (.D(n9[3]), .SP(sys_clk_enable_236), 
            .CD(n40166), .CK(sys_clk), .Q(tx_byte_index[3]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam tx_byte_index_6622__i3.GSR = "ENABLED";
    FD1P3IX tx_byte_index_6622__i2 (.D(n9[2]), .SP(sys_clk_enable_236), 
            .CD(n40166), .CK(sys_clk), .Q(tx_byte_index[2]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam tx_byte_index_6622__i2.GSR = "ENABLED";
    FD1P3IX tx_byte_index_6622__i1 (.D(n9[1]), .SP(sys_clk_enable_236), 
            .CD(n40166), .CK(sys_clk), .Q(\tx_byte_index[1] ));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam tx_byte_index_6622__i1.GSR = "ENABLED";
    FD1P3IX tx_word_index_6624__i0 (.D(n8[0]), .SP(sys_clk_enable_217), 
            .CD(n40212), .CK(sys_clk), .Q(tx_word_index[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(371[42:62])
    defparam tx_word_index_6624__i0.GSR = "ENABLED";
    PFUMX i40075 (.BLUT(n50859), .ALUT(n50858), .C0(\tx_byte_index[0] ), 
          .Z(n50860));
    FD1P3IX dat_i_i1 (.D(n48589), .SP(sys_clk_enable_246), .CD(n38023), 
            .CK(sys_clk), .Q(dat_i[1])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=64, LSE_RCOL=6, LSE_LLINE=528, LSE_RLINE=562 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam dat_i_i1.GSR = "ENABLED";
    FD1P3AX dat_i_i2 (.D(next_dat_i_15__N_4452[2]), .SP(sys_clk_enable_246), 
            .CK(sys_clk), .Q(dat_i[2])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=64, LSE_RCOL=6, LSE_LLINE=528, LSE_RLINE=562 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam dat_i_i2.GSR = "ENABLED";
    FD1P3AX dat_i_i3 (.D(\next_dat_i_15__N_4452[3] ), .SP(sys_clk_enable_246), 
            .CK(sys_clk), .Q(dat_i[3])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=64, LSE_RCOL=6, LSE_LLINE=528, LSE_RLINE=562 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam dat_i_i3.GSR = "ENABLED";
    FD1P3AX dat_i_i6 (.D(next_dat_i_15__N_4452[6]), .SP(sys_clk_enable_246), 
            .CK(sys_clk), .Q(dat_i[6])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=64, LSE_RCOL=6, LSE_LLINE=528, LSE_RLINE=562 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam dat_i_i6.GSR = "ENABLED";
    FD1P3IX tx_byte_index_6622__i0 (.D(n52395), .SP(sys_clk_enable_236), 
            .CD(n40166), .CK(sys_clk), .Q(\tx_byte_index[0] ));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(327[42:62])
    defparam tx_byte_index_6622__i0.GSR = "ENABLED";
    FD1P3IX dat_i_i0 (.D(n48731), .SP(sys_clk_enable_246), .CD(n38023), 
            .CK(sys_clk), .Q(dat_i[0])) /* synthesis LSE_LINE_FILE_ID=6, LSE_LCOL=64, LSE_RCOL=6, LSE_LLINE=528, LSE_RLINE=562 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(198[14] 210[12])
    defparam dat_i_i0.GSR = "ENABLED";
    \uart_core(CLK_IN_MHZ=38)  uart_core_inst (.sys_clk(sys_clk), .\next_state_9__N_4551[6] (next_state_9__N_4551[6]), 
            .\next_state_4__N_1567[2] (\next_state_4__N_1567[2] ), .\next_state_9__N_4531[5] (next_state_9__N_4531[5]), 
            .GND_net(GND_net), .sout_c(sout_c), .n22616(n22616), .n38171(n38171), 
            .n36607(n36607), .\next_state_9__N_4478[7] (next_state_9__N_4478[7]), 
            .sin_c(sin_c), .n53885(n53885), .\adr_i[0] (adr_i[0]), .cyc_i(cyc_i), 
            .we_i(we_i), .\adr_i[1] (adr_i[1]), .\adr_i[2] (adr_i[2]), 
            .\dat_i[0] (dat_i[0]), .\next_state_9__N_4541[6] (next_state_9__N_4541[6]), 
            .rxrdy_n_c(rxrdy_n_c), .\dat_i[1] (dat_i[1]), .\dat_i[2] (dat_i[2]), 
            .\dat_i[3] (dat_i[3]), .\dat_i[5] (dat_i[5]), .\dat_i[6] (dat_i[6]), 
            .n53884(n53884)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_top.v(114[5] 160[6])
    
endmodule
//
// Verilog Description of module \uart_core(CLK_IN_MHZ=38) 
//

module \uart_core(CLK_IN_MHZ=38)  (sys_clk, \next_state_9__N_4551[6] , \next_state_4__N_1567[2] , 
            \next_state_9__N_4531[5] , GND_net, sout_c, n22616, n38171, 
            n36607, \next_state_9__N_4478[7] , sin_c, n53885, \adr_i[0] , 
            cyc_i, we_i, \adr_i[1] , \adr_i[2] , \dat_i[0] , \next_state_9__N_4541[6] , 
            rxrdy_n_c, \dat_i[1] , \dat_i[2] , \dat_i[3] , \dat_i[5] , 
            \dat_i[6] , n53884) /* synthesis syn_module_defined=1 */ ;
    input sys_clk;
    output \next_state_9__N_4551[6] ;
    input \next_state_4__N_1567[2] ;
    output \next_state_9__N_4531[5] ;
    input GND_net;
    output sout_c;
    input n22616;
    input n38171;
    input n36607;
    output \next_state_9__N_4478[7] ;
    input sin_c;
    input n53885;
    input \adr_i[0] ;
    input cyc_i;
    input we_i;
    input \adr_i[1] ;
    input \adr_i[2] ;
    input \dat_i[0] ;
    output \next_state_9__N_4541[6] ;
    output rxrdy_n_c;
    input \dat_i[1] ;
    input \dat_i[2] ;
    input \dat_i[3] ;
    input \dat_i[5] ;
    input \dat_i[6] ;
    input n53884;
    
    wire sys_clk /* synthesis SET_AS_NETWORK=sys_clk, is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(220[10:17])
    wire [15:0]divisor;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_core.v(158[23:30])
    wire [6:0]lcr;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/intface.v(172[15:18])
    wire [1:0]databits;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_core.v(136[23:31])
    wire [6:0]n15;
    wire [7:0]THR;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_core.v(135[23:26])
    
    wire thr_wr, rx_rdy, rbr_rd;
    
    \txmitt(DATAWIDTH=8)  u_txmitt (.\divisor[8] (divisor[8]), .\divisor[4] (divisor[4]), 
            .\divisor[6] (divisor[6]), .\divisor[3] (divisor[3]), .\divisor[2] (divisor[2]), 
            .\divisor[1] (divisor[1]), .\divisor[0] (divisor[0]), .sys_clk(sys_clk), 
            .\lcr[2] (lcr[2]), .databits({databits}), .parity_en(n15[3]), 
            .\next_state_9__N_4551[6] (\next_state_9__N_4551[6] ), .\next_state_4__N_1567[2] (\next_state_4__N_1567[2] ), 
            .\next_state_9__N_4531[5] (\next_state_9__N_4531[5] ), .GND_net(GND_net), 
            .tx_break(n15[6]), .sout_c(sout_c), .\THR[1] (THR[1]), .\THR[2] (THR[2]), 
            .\THR[3] (THR[3]), .\THR[4] (THR[4]), .\THR[6] (THR[6]), .\THR[0] (THR[0]), 
            .parity_even(n15[4]), .thr_wr(thr_wr), .n22616(n22616), .n38171(n38171), 
            .n36607(n36607), .\next_state_9__N_4478[7] (\next_state_9__N_4478[7] )) /* synthesis syn_module_defined=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_core.v(283[7] 300[4])
    \rxcver(FIFO=0)  u_rxcver (.parity_en(n15[3]), .sys_clk(sys_clk), .sin_c(sin_c), 
            .rx_rdy(rx_rdy), .rbr_rd(rbr_rd), .n53885(n53885), .databits({databits}), 
            .GND_net(GND_net), .\divisor[8] (divisor[8]), .\divisor[4] (divisor[4]), 
            .\divisor[6] (divisor[6]), .\divisor[3] (divisor[3]), .\divisor[1] (divisor[1]), 
            .\divisor[2] (divisor[2]), .\divisor[0] (divisor[0])) /* synthesis syn_module_defined=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_core.v(259[6] 279[4])
    \intface(CLK_IN_MHZ=38)  u_intface (.\adr_i[0] (\adr_i[0] ), .cyc_i(cyc_i), 
            .we_i(we_i), .\adr_i[1] (\adr_i[1] ), .\adr_i[2] (\adr_i[2] ), 
            .\THR[0] (THR[0]), .sys_clk(sys_clk), .\dat_i[0] (\dat_i[0] ), 
            .databits({databits}), .\divisor[0] (divisor[0]), .thr_wr(thr_wr), 
            .rbr_rd(rbr_rd), .\next_state_9__N_4541[6] (\next_state_9__N_4541[6] ), 
            .n53885(n53885), .rx_rdy(rx_rdy), .rxrdy_n_c(rxrdy_n_c), .\THR[1] (THR[1]), 
            .\dat_i[1] (\dat_i[1] ), .\THR[2] (THR[2]), .\dat_i[2] (\dat_i[2] ), 
            .\THR[3] (THR[3]), .\dat_i[3] (\dat_i[3] ), .\THR[4] (THR[4]), 
            .\dat_i[5] (\dat_i[5] ), .\THR[6] (THR[6]), .\dat_i[6] (\dat_i[6] ), 
            .\lcr[2] (lcr[2]), .parity_en(n15[3]), .parity_even(n15[4]), 
            .tx_break(n15[6]), .\divisor[1] (divisor[1]), .\divisor[2] (divisor[2]), 
            .\divisor[3] (divisor[3]), .\divisor[4] (divisor[4]), .\divisor[6] (divisor[6]), 
            .\divisor[8] (divisor[8]), .n53884(n53884)) /* synthesis syn_module_defined=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_core.v(169[10] 209[4])
    
endmodule
//
// Verilog Description of module \txmitt(DATAWIDTH=8) 
//

module \txmitt(DATAWIDTH=8)  (\divisor[8] , \divisor[4] , \divisor[6] , 
            \divisor[3] , \divisor[2] , \divisor[1] , \divisor[0] , 
            sys_clk, \lcr[2] , databits, parity_en, \next_state_9__N_4551[6] , 
            \next_state_4__N_1567[2] , \next_state_9__N_4531[5] , GND_net, 
            tx_break, sout_c, \THR[1] , \THR[2] , \THR[3] , \THR[4] , 
            \THR[6] , \THR[0] , parity_even, thr_wr, n22616, n38171, 
            n36607, \next_state_9__N_4478[7] ) /* synthesis syn_module_defined=1 */ ;
    input \divisor[8] ;
    input \divisor[4] ;
    input \divisor[6] ;
    input \divisor[3] ;
    input \divisor[2] ;
    input \divisor[1] ;
    input \divisor[0] ;
    input sys_clk;
    input \lcr[2] ;
    input [1:0]databits;
    input parity_en;
    output \next_state_9__N_4551[6] ;
    input \next_state_4__N_1567[2] ;
    output \next_state_9__N_4531[5] ;
    input GND_net;
    input tx_break;
    output sout_c;
    input \THR[1] ;
    input \THR[2] ;
    input \THR[3] ;
    input \THR[4] ;
    input \THR[6] ;
    input \THR[0] ;
    input parity_even;
    input thr_wr;
    input n22616;
    input n38171;
    input n36607;
    output \next_state_9__N_4478[7] ;
    
    wire sys_clk /* synthesis SET_AS_NETWORK=sys_clk, is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(220[10:17])
    wire [2:0]tx_cnt;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(102[28:34])
    wire [15:0]counter;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(118[14:21])
    
    wire n47341;
    wire [2:0]tx_cnt_2__N_5022;
    
    wire n52202;
    wire [2:0]tx_state;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(117[13:21])
    
    wire n21, sys_clk_enable_239, n6, n48115, n11;
    wire [15:0]n1;
    
    wire n52544, n52408, n52543, n52547, n52187, n52546, n52550, 
        n52549, n52553, n52552, n52556, n52555, n52559, n52558, 
        n52589, n52588, sys_clk_enable_237, n52560, n52601, n52600, 
        n52604, n52603;
    wire [7:0]tsr;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(91[28:31])
    
    wire sys_clk_enable_135;
    wire [7:0]tsr_7__N_4939;
    
    wire tx_parity, tx_parity_N_5052, tx_in_shift_s1, tx_in_shift_s, 
        tx_in_shift_s_N_5066, n16225, n43877, n43876, n5, n43875, 
        tx_output, n43874, n43873, n43872, n43871, n30763, n43870, 
        n14_adj_5100, n12, tx_output_N_5048, n52186, n28_adj_5101, 
        n24_adj_5102, n16_adj_5103, n26_adj_5104, n20_adj_5105, n52605;
    wire [2:0]tx_state_2__N_4950;
    
    wire n46457, n52557, n52554, n52551, n52548, n52590, n52545, 
        n52602, sys_clk_enable_238;
    
    LUT4 i33228_4_lut_4_lut (.A(tx_cnt[0]), .B(tx_cnt[1]), .C(counter[0]), 
         .D(n47341), .Z(tx_cnt_2__N_5022[1])) /* synthesis lut_function=(A (B ((D)+!C)+!B !((D)+!C))+!A (B)) */ ;
    defparam i33228_4_lut_4_lut.init = 16'hcc6c;
    LUT4 i1_4_lut_4_lut (.A(n52202), .B(tx_state[1]), .C(n21), .D(tx_state[2]), 
         .Z(sys_clk_enable_239)) /* synthesis lut_function=(A (C)+!A (B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam i1_4_lut_4_lut.init = 16'hf5f4;
    LUT4 i33226_4_lut_4_lut (.A(n52202), .B(tx_cnt[0]), .C(tx_cnt[1]), 
         .D(tx_cnt[2]), .Z(tx_cnt_2__N_5022[2])) /* synthesis lut_function=(A (D)+!A !(B (C (D)+!C !(D))+!B !(D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam i33226_4_lut_4_lut.init = 16'hbf40;
    LUT4 i1_4_lut_4_lut_adj_144 (.A(n52202), .B(tx_cnt[2]), .C(n6), .D(n48115), 
         .Z(n11)) /* synthesis lut_function=(A (D)+!A (B (C+(D))+!B (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam i1_4_lut_4_lut_adj_144.init = 16'hff40;
    LUT4 mux_3398_i8_then_1_lut (.A(n1[7]), .Z(n52544)) /* synthesis lut_function=(A) */ ;
    defparam mux_3398_i8_then_1_lut.init = 16'haaaa;
    LUT4 mux_3398_i8_else_1_lut (.A(tx_state[2]), .B(counter[0]), .C(n52408), 
         .D(\divisor[8] ), .Z(n52543)) /* synthesis lut_function=(!((B+!(C (D)))+!A)) */ ;
    defparam mux_3398_i8_else_1_lut.init = 16'h2000;
    LUT4 mux_3398_i6_then_1_lut (.A(n1[5]), .Z(n52547)) /* synthesis lut_function=(A) */ ;
    defparam mux_3398_i6_then_1_lut.init = 16'haaaa;
    LUT4 mux_3398_i6_else_1_lut (.A(\divisor[4] ), .B(counter[0]), .C(\divisor[6] ), 
         .D(n52187), .Z(n52546)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;
    defparam mux_3398_i6_else_1_lut.init = 16'h3022;
    LUT4 mux_3398_i4_then_1_lut (.A(n1[3]), .Z(n52550)) /* synthesis lut_function=(A) */ ;
    defparam mux_3398_i4_then_1_lut.init = 16'haaaa;
    LUT4 mux_3398_i4_else_1_lut (.A(\divisor[3] ), .B(counter[0]), .C(\divisor[4] ), 
         .D(n52187), .Z(n52549)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;
    defparam mux_3398_i4_else_1_lut.init = 16'h3022;
    LUT4 mux_3398_i3_then_1_lut (.A(n1[2]), .Z(n52553)) /* synthesis lut_function=(A) */ ;
    defparam mux_3398_i3_then_1_lut.init = 16'haaaa;
    LUT4 mux_3398_i3_else_1_lut (.A(\divisor[2] ), .B(counter[0]), .C(\divisor[3] ), 
         .D(n52187), .Z(n52552)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;
    defparam mux_3398_i3_else_1_lut.init = 16'h3022;
    LUT4 mux_3398_i2_then_1_lut (.A(n1[1]), .Z(n52556)) /* synthesis lut_function=(A) */ ;
    defparam mux_3398_i2_then_1_lut.init = 16'haaaa;
    LUT4 mux_3398_i2_else_1_lut (.A(\divisor[1] ), .B(counter[0]), .C(\divisor[2] ), 
         .D(n52187), .Z(n52555)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;
    defparam mux_3398_i2_else_1_lut.init = 16'h3022;
    LUT4 mux_3398_i1_then_1_lut (.A(n1[0]), .Z(n52559)) /* synthesis lut_function=(A) */ ;
    defparam mux_3398_i1_then_1_lut.init = 16'haaaa;
    LUT4 mux_3398_i1_else_1_lut (.A(\divisor[0] ), .B(counter[0]), .C(\divisor[1] ), 
         .D(n52187), .Z(n52558)) /* synthesis lut_function=(!(A (B+!(C+!(D)))+!A (B+!(C (D))))) */ ;
    defparam mux_3398_i1_else_1_lut.init = 16'h3022;
    LUT4 i40577_then_1_lut (.A(n1[6]), .Z(n52589)) /* synthesis lut_function=(A) */ ;
    defparam i40577_then_1_lut.init = 16'haaaa;
    LUT4 i40577_else_1_lut (.A(tx_state[2]), .B(counter[0]), .C(n52408), 
         .D(\divisor[6] ), .Z(n52588)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A (B+!(D)))) */ ;
    defparam i40577_else_1_lut.init = 16'h1300;
    FD1P3AX counter_i0_i0 (.D(n52560), .SP(sys_clk_enable_237), .CK(sys_clk), 
            .Q(counter[0])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=7, LSE_RCOL=4, LSE_LLINE=283, LSE_RLINE=300 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam counter_i0_i0.GSR = "ENABLED";
    LUT4 i40574_then_1_lut (.A(n1[8]), .Z(n52601)) /* synthesis lut_function=(A) */ ;
    defparam i40574_then_1_lut.init = 16'haaaa;
    LUT4 i40574_else_1_lut (.A(tx_state[2]), .B(counter[0]), .C(n52408), 
         .D(\divisor[8] ), .Z(n52600)) /* synthesis lut_function=(!(A (B+(C+!(D)))+!A (B+!(D)))) */ ;
    defparam i40574_else_1_lut.init = 16'h1300;
    LUT4 lcr_2__bdd_4_lut_then_3_lut (.A(\lcr[2] ), .B(databits[0]), .C(databits[1]), 
         .Z(n52604)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;
    defparam lcr_2__bdd_4_lut_then_3_lut.init = 16'h0202;
    LUT4 lcr_2__bdd_4_lut_else_3_lut (.A(tx_state[0]), .B(parity_en), .Z(n52603)) /* synthesis lut_function=(!((B)+!A)) */ ;
    defparam lcr_2__bdd_4_lut_else_3_lut.init = 16'h2222;
    FD1P3AX tsr_i0 (.D(tsr_7__N_4939[0]), .SP(sys_clk_enable_135), .CK(sys_clk), 
            .Q(tsr[0])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=7, LSE_RCOL=4, LSE_LLINE=283, LSE_RLINE=300 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam tsr_i0.GSR = "ENABLED";
    FD1P3AY tx_parity_129 (.D(tx_parity_N_5052), .SP(sys_clk_enable_135), 
            .CK(sys_clk), .Q(tx_parity)) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=7, LSE_RCOL=4, LSE_LLINE=283, LSE_RLINE=300 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam tx_parity_129.GSR = "ENABLED";
    FD1S3AX tx_in_shift_s1_134 (.D(tx_in_shift_s), .CK(sys_clk), .Q(tx_in_shift_s1)) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=7, LSE_RCOL=4, LSE_LLINE=283, LSE_RLINE=300 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(472[14] 475[14])
    defparam tx_in_shift_s1_134.GSR = "ENABLED";
    FD1S3AX tx_in_shift_s_136 (.D(tx_in_shift_s_N_5066), .CK(sys_clk), .Q(tx_in_shift_s)) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=7, LSE_RCOL=4, LSE_LLINE=283, LSE_RLINE=300 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(486[14] 489[33])
    defparam tx_in_shift_s_136.GSR = "ENABLED";
    LUT4 i1_2_lut (.A(\next_state_9__N_4551[6] ), .B(\next_state_4__N_1567[2] ), 
         .Z(\next_state_9__N_4531[5] )) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(452[11] 455[26])
    defparam i1_2_lut.init = 16'h8888;
    FD1S3AY thr_empty_133 (.D(n16225), .CK(sys_clk), .Q(\next_state_9__N_4551[6] )) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=7, LSE_RCOL=4, LSE_LLINE=283, LSE_RLINE=300 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(452[11] 455[26])
    defparam thr_empty_133.GSR = "ENABLED";
    CCU2D sub_10_add_2_17 (.A0(counter[15]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n43877), .S0(n1[15]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(304[24:38])
    defparam sub_10_add_2_17.INIT0 = 16'h5555;
    defparam sub_10_add_2_17.INIT1 = 16'h0000;
    defparam sub_10_add_2_17.INJECT1_0 = "NO";
    defparam sub_10_add_2_17.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_15 (.A0(counter[13]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(counter[14]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43876), .COUT(n43877), .S0(n1[13]), .S1(n1[14]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(304[24:38])
    defparam sub_10_add_2_15.INIT0 = 16'h5555;
    defparam sub_10_add_2_15.INIT1 = 16'h5555;
    defparam sub_10_add_2_15.INJECT1_0 = "NO";
    defparam sub_10_add_2_15.INJECT1_1 = "NO";
    LUT4 i37681_3_lut (.A(tx_state[2]), .B(tx_state[1]), .C(\next_state_9__N_4551[6] ), 
         .Z(n5)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam i37681_3_lut.init = 16'h0101;
    CCU2D sub_10_add_2_13 (.A0(counter[11]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(counter[12]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43875), .COUT(n43876), .S0(n1[11]), .S1(n1[12]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(304[24:38])
    defparam sub_10_add_2_13.INIT0 = 16'h5555;
    defparam sub_10_add_2_13.INIT1 = 16'h5555;
    defparam sub_10_add_2_13.INJECT1_0 = "NO";
    defparam sub_10_add_2_13.INJECT1_1 = "NO";
    LUT4 i25903_2_lut (.A(tx_output), .B(tx_break), .Z(sout_c)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(515[16:51])
    defparam i25903_2_lut.init = 16'h2222;
    CCU2D sub_10_add_2_11 (.A0(counter[9]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(counter[10]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43874), .COUT(n43875), .S0(n1[9]), .S1(n1[10]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(304[24:38])
    defparam sub_10_add_2_11.INIT0 = 16'h5555;
    defparam sub_10_add_2_11.INIT1 = 16'h5555;
    defparam sub_10_add_2_11.INJECT1_0 = "NO";
    defparam sub_10_add_2_11.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_9 (.A0(counter[7]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(counter[8]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43873), .COUT(n43874), .S0(n1[7]), .S1(n1[8]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(304[24:38])
    defparam sub_10_add_2_9.INIT0 = 16'h5555;
    defparam sub_10_add_2_9.INIT1 = 16'h5555;
    defparam sub_10_add_2_9.INJECT1_0 = "NO";
    defparam sub_10_add_2_9.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_7 (.A0(counter[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(counter[6]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43872), .COUT(n43873), .S0(n1[5]), .S1(n1[6]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(304[24:38])
    defparam sub_10_add_2_7.INIT0 = 16'h5555;
    defparam sub_10_add_2_7.INIT1 = 16'h5555;
    defparam sub_10_add_2_7.INJECT1_0 = "NO";
    defparam sub_10_add_2_7.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_5 (.A0(counter[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(counter[4]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43871), .COUT(n43872), .S0(n1[3]), .S1(n1[4]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(304[24:38])
    defparam sub_10_add_2_5.INIT0 = 16'h5555;
    defparam sub_10_add_2_5.INIT1 = 16'h5555;
    defparam sub_10_add_2_5.INJECT1_0 = "NO";
    defparam sub_10_add_2_5.INJECT1_1 = "NO";
    LUT4 tx_state_1__bdd_3_lut_rep_379 (.A(tx_state[1]), .B(tx_state[2]), 
         .C(tx_state[0]), .Z(sys_clk_enable_237)) /* synthesis lut_function=(!(A (B (C))+!A !(B+(C)))) */ ;
    defparam tx_state_1__bdd_3_lut_rep_379.init = 16'h7e7e;
    LUT4 i20092_2_lut_4_lut (.A(tx_state[1]), .B(tx_state[2]), .C(tx_state[0]), 
         .D(n47341), .Z(n30763)) /* synthesis lut_function=(!(A (B (C+(D))+!B (D))+!A (B (D)+!B ((D)+!C)))) */ ;
    defparam i20092_2_lut_4_lut.init = 16'h007e;
    CCU2D sub_10_add_2_3 (.A0(counter[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(counter[2]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43870), .COUT(n43871), .S0(n1[1]), .S1(n1[2]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(304[24:38])
    defparam sub_10_add_2_3.INIT0 = 16'h5555;
    defparam sub_10_add_2_3.INIT1 = 16'h5555;
    defparam sub_10_add_2_3.INJECT1_0 = "NO";
    defparam sub_10_add_2_3.INJECT1_1 = "NO";
    CCU2D sub_10_add_2_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), .D0(GND_net), 
          .A1(counter[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n43870), .S1(n1[0]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(304[24:38])
    defparam sub_10_add_2_1.INIT0 = 16'hF000;
    defparam sub_10_add_2_1.INIT1 = 16'h5555;
    defparam sub_10_add_2_1.INJECT1_0 = "NO";
    defparam sub_10_add_2_1.INJECT1_1 = "NO";
    LUT4 i2_3_lut_rep_251_4_lut (.A(counter[0]), .B(n47341), .C(n52408), 
         .D(tx_state[2]), .Z(n52187)) /* synthesis lut_function=(!(A+(B+!(C (D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam i2_3_lut_rep_251_4_lut.init = 16'h1000;
    LUT4 i19022_3_lut (.A(tsr[2]), .B(\THR[1] ), .C(tx_state[2]), .Z(tsr_7__N_4939[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(287[9] 392[16])
    defparam i19022_3_lut.init = 16'hcaca;
    LUT4 i19020_3_lut (.A(tsr[3]), .B(\THR[2] ), .C(tx_state[2]), .Z(tsr_7__N_4939[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(287[9] 392[16])
    defparam i19020_3_lut.init = 16'hcaca;
    LUT4 i19018_3_lut (.A(tsr[4]), .B(\THR[3] ), .C(tx_state[2]), .Z(tsr_7__N_4939[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(287[9] 392[16])
    defparam i19018_3_lut.init = 16'hcaca;
    LUT4 i19016_3_lut (.A(tsr[5]), .B(\THR[4] ), .C(tx_state[2]), .Z(tsr_7__N_4939[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(287[9] 392[16])
    defparam i19016_3_lut.init = 16'hcaca;
    LUT4 i19014_3_lut (.A(tsr[6]), .B(\THR[4] ), .C(tx_state[2]), .Z(tsr_7__N_4939[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(287[9] 392[16])
    defparam i19014_3_lut.init = 16'hcaca;
    PFUMX i26 (.BLUT(n14_adj_5100), .ALUT(n12), .C0(tx_state[1]), .Z(tx_output_N_5048));
    LUT4 i27195_2_lut (.A(\THR[6] ), .B(tx_state[2]), .Z(tsr_7__N_4939[6])) /* synthesis lut_function=(A (B)) */ ;
    defparam i27195_2_lut.init = 16'h8888;
    LUT4 i2_3_lut_rep_250_4_lut (.A(counter[0]), .B(n47341), .C(tx_state[0]), 
         .D(n48115), .Z(n52186)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam i2_3_lut_rep_250_4_lut.init = 16'h0200;
    LUT4 i2_4_lut (.A(databits[1]), .B(databits[0]), .C(tx_cnt[1]), .D(tx_cnt[0]), 
         .Z(n6)) /* synthesis lut_function=(A (B (C (D))+!B !((D)+!C))+!A !(B (C+!(D))+!B (C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(117[13:21])
    defparam i2_4_lut.init = 16'h8421;
    LUT4 i1_4_lut (.A(tx_state[2]), .B(n52186), .C(n52202), .D(n52408), 
         .Z(sys_clk_enable_135)) /* synthesis lut_function=(A (B)+!A (B+!(C+!(D)))) */ ;
    defparam i1_4_lut.init = 16'hcdcc;
    LUT4 i19009_3_lut (.A(tsr[1]), .B(\THR[0] ), .C(tx_state[2]), .Z(tsr_7__N_4939[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(287[9] 392[16])
    defparam i19009_3_lut.init = 16'hcaca;
    LUT4 i1_2_lut_adj_145 (.A(tx_state[2]), .B(tx_state[1]), .Z(n48115)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(117[13:21])
    defparam i1_2_lut_adj_145.init = 16'h8888;
    LUT4 i14_4_lut (.A(counter[1]), .B(n28_adj_5101), .C(n24_adj_5102), 
         .D(n16_adj_5103), .Z(n47341)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam i14_4_lut.init = 16'hfffe;
    LUT4 i13_4_lut (.A(counter[11]), .B(n26_adj_5104), .C(n20_adj_5105), 
         .D(counter[6]), .Z(n28_adj_5101)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam i13_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_rep_472 (.A(tx_state[0]), .B(tx_state[1]), .Z(n52408)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam i1_2_lut_rep_472.init = 16'h2222;
    LUT4 i1_2_lut_3_lut (.A(tx_state[0]), .B(tx_state[1]), .C(tx_state[2]), 
         .Z(tx_in_shift_s_N_5066)) /* synthesis lut_function=(!((B+(C))+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam i1_2_lut_3_lut.init = 16'h0202;
    LUT4 i9_4_lut (.A(counter[14]), .B(counter[15]), .C(counter[4]), .D(counter[2]), 
         .Z(n24_adj_5102)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam i9_4_lut.init = 16'hfffe;
    LUT4 i1_2_lut_adj_146 (.A(counter[13]), .B(counter[5]), .Z(n16_adj_5103)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam i1_2_lut_adj_146.init = 16'heeee;
    LUT4 i1_3_lut_3_lut_4_lut (.A(tx_state[0]), .B(tx_state[1]), .C(n52605), 
         .D(tx_state[2]), .Z(tx_state_2__N_4950[0])) /* synthesis lut_function=(!(A ((D)+!C)+!A !(B+!((D)+!C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(287[9] 392[16])
    defparam i1_3_lut_3_lut_4_lut.init = 16'h44f4;
    LUT4 i11_4_lut (.A(counter[7]), .B(counter[3]), .C(counter[10]), .D(counter[8]), 
         .Z(n26_adj_5104)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam i11_4_lut.init = 16'hfffe;
    LUT4 i5_2_lut (.A(counter[12]), .B(counter[9]), .Z(n20_adj_5105)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam i5_2_lut.init = 16'heeee;
    LUT4 i19007_4_lut (.A(tx_parity), .B(parity_even), .C(tx_state[2]), 
         .D(tsr[0]), .Z(tx_parity_N_5052)) /* synthesis lut_function=(!(A (B (C+(D))+!B !(C+!(D)))+!A (B (C+!(D))+!B !(C+(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(287[9] 392[16])
    defparam i19007_4_lut.init = 16'h353a;
    LUT4 i25758_4_lut (.A(\next_state_9__N_4551[6] ), .B(thr_wr), .C(tx_in_shift_s), 
         .D(tx_in_shift_s1), .Z(n16225)) /* synthesis lut_function=(!(A (B)+!A (B+((D)+!C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(452[11] 455[26])
    defparam i25758_4_lut.init = 16'h2232;
    LUT4 i11_4_lut_4_lut (.A(\divisor[4] ), .B(counter[0]), .C(n47341), 
         .D(n1[4]), .Z(n46457)) /* synthesis lut_function=(A (B (C (D))+!B ((D)+!C))+!A (C (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(287[9] 392[16])
    defparam i11_4_lut_4_lut.init = 16'hf202;
    FD1P3AX counter_i0_i1 (.D(n52557), .SP(sys_clk_enable_237), .CK(sys_clk), 
            .Q(counter[1])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=7, LSE_RCOL=4, LSE_LLINE=283, LSE_RLINE=300 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam counter_i0_i1.GSR = "ENABLED";
    LUT4 i39943_3_lut (.A(tx_state[2]), .B(tx_state[1]), .C(tx_state[0]), 
         .Z(tx_state_2__N_4950[1])) /* synthesis lut_function=(!(A+(B (C)))) */ ;
    defparam i39943_3_lut.init = 16'h1515;
    LUT4 i1_4_lut_4_lut_adj_147 (.A(tx_state[2]), .B(tx_state[1]), .C(\lcr[2] ), 
         .D(tx_state[0]), .Z(tx_state_2__N_4950[2])) /* synthesis lut_function=(!(A+!(B (C (D))+!B !(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(287[9] 392[16])
    defparam i1_4_lut_4_lut_adj_147.init = 16'h4011;
    LUT4 i1_4_lut_4_lut_4_lut (.A(tx_state[2]), .B(tx_state[0]), .C(tx_parity), 
         .D(parity_even), .Z(n12)) /* synthesis lut_function=(!(A+!(B+!((D)+!C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(287[9] 392[16])
    defparam i1_4_lut_4_lut_4_lut.init = 16'h4454;
    FD1P3AX counter_i0_i2 (.D(n52554), .SP(sys_clk_enable_237), .CK(sys_clk), 
            .Q(counter[2])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=7, LSE_RCOL=4, LSE_LLINE=283, LSE_RLINE=300 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam counter_i0_i2.GSR = "ENABLED";
    FD1P3AX counter_i0_i3 (.D(n52551), .SP(sys_clk_enable_237), .CK(sys_clk), 
            .Q(counter[3])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=7, LSE_RCOL=4, LSE_LLINE=283, LSE_RLINE=300 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam counter_i0_i3.GSR = "ENABLED";
    FD1P3AX counter_i0_i4 (.D(n46457), .SP(sys_clk_enable_237), .CK(sys_clk), 
            .Q(counter[4])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=7, LSE_RCOL=4, LSE_LLINE=283, LSE_RLINE=300 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam counter_i0_i4.GSR = "ENABLED";
    FD1P3AX counter_i0_i5 (.D(n52548), .SP(sys_clk_enable_237), .CK(sys_clk), 
            .Q(counter[5])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=7, LSE_RCOL=4, LSE_LLINE=283, LSE_RLINE=300 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam counter_i0_i5.GSR = "ENABLED";
    FD1P3AX counter_i0_i6 (.D(n52590), .SP(sys_clk_enable_237), .CK(sys_clk), 
            .Q(counter[6])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=7, LSE_RCOL=4, LSE_LLINE=283, LSE_RLINE=300 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam counter_i0_i6.GSR = "ENABLED";
    FD1P3AX counter_i0_i7 (.D(n52545), .SP(sys_clk_enable_237), .CK(sys_clk), 
            .Q(counter[7])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=7, LSE_RCOL=4, LSE_LLINE=283, LSE_RLINE=300 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam counter_i0_i7.GSR = "ENABLED";
    FD1P3AX counter_i0_i8 (.D(n52602), .SP(sys_clk_enable_237), .CK(sys_clk), 
            .Q(counter[8])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=7, LSE_RCOL=4, LSE_LLINE=283, LSE_RLINE=300 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam counter_i0_i8.GSR = "ENABLED";
    FD1P3AX tsr_i1 (.D(tsr_7__N_4939[1]), .SP(sys_clk_enable_135), .CK(sys_clk), 
            .Q(tsr[1])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=7, LSE_RCOL=4, LSE_LLINE=283, LSE_RLINE=300 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam tsr_i1.GSR = "ENABLED";
    FD1P3AX tsr_i2 (.D(tsr_7__N_4939[2]), .SP(sys_clk_enable_135), .CK(sys_clk), 
            .Q(tsr[2])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=7, LSE_RCOL=4, LSE_LLINE=283, LSE_RLINE=300 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam tsr_i2.GSR = "ENABLED";
    FD1P3AX tsr_i3 (.D(tsr_7__N_4939[3]), .SP(sys_clk_enable_135), .CK(sys_clk), 
            .Q(tsr[3])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=7, LSE_RCOL=4, LSE_LLINE=283, LSE_RLINE=300 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam tsr_i3.GSR = "ENABLED";
    FD1P3AX tsr_i4 (.D(tsr_7__N_4939[4]), .SP(sys_clk_enable_135), .CK(sys_clk), 
            .Q(tsr[4])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=7, LSE_RCOL=4, LSE_LLINE=283, LSE_RLINE=300 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam tsr_i4.GSR = "ENABLED";
    FD1P3AX tsr_i5 (.D(tsr_7__N_4939[5]), .SP(sys_clk_enable_135), .CK(sys_clk), 
            .Q(tsr[5])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=7, LSE_RCOL=4, LSE_LLINE=283, LSE_RLINE=300 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam tsr_i5.GSR = "ENABLED";
    FD1P3AX tsr_i6 (.D(tsr_7__N_4939[6]), .SP(sys_clk_enable_135), .CK(sys_clk), 
            .Q(tsr[6])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=7, LSE_RCOL=4, LSE_LLINE=283, LSE_RLINE=300 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam tsr_i6.GSR = "ENABLED";
    LUT4 i1_2_lut_adj_148 (.A(tx_state[2]), .B(tsr[0]), .Z(n14_adj_5100)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(287[9] 392[16])
    defparam i1_2_lut_adj_148.init = 16'heeee;
    LUT4 i1_2_lut_rep_266 (.A(counter[0]), .B(n47341), .Z(n52202)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam i1_2_lut_rep_266.init = 16'hdddd;
    PFUMX i27 (.BLUT(n5), .ALUT(n11), .C0(tx_state[0]), .Z(n21));
    LUT4 i3_4_lut (.A(\next_state_9__N_4551[6] ), .B(n22616), .C(n38171), 
         .D(n36607), .Z(\next_state_9__N_4478[7] )) /* synthesis lut_function=(!(A+((C+(D))+!B))) */ ;
    defparam i3_4_lut.init = 16'h0004;
    LUT4 i30271_3_lut_4_lut_3_lut (.A(counter[0]), .B(n47341), .C(tx_cnt[0]), 
         .Z(tx_cnt_2__N_5022[0])) /* synthesis lut_function=(A (B (C)+!B !(C))+!A (C)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam i30271_3_lut_4_lut_3_lut.init = 16'hd2d2;
    LUT4 i1_2_lut_4_lut (.A(n52202), .B(n48115), .C(tx_state[0]), .D(tx_in_shift_s_N_5066), 
         .Z(sys_clk_enable_238)) /* synthesis lut_function=(A (D)+!A (B ((D)+!C)+!B (D))) */ ;
    defparam i1_2_lut_4_lut.init = 16'hff04;
    PFUMX i40996 (.BLUT(n52603), .ALUT(n52604), .C0(tx_state[1]), .Z(n52605));
    PFUMX i40994 (.BLUT(n52600), .ALUT(n52601), .C0(n47341), .Z(n52602));
    PFUMX i40986 (.BLUT(n52588), .ALUT(n52589), .C0(n47341), .Z(n52590));
    PFUMX i40966 (.BLUT(n52558), .ALUT(n52559), .C0(n47341), .Z(n52560));
    PFUMX i40964 (.BLUT(n52555), .ALUT(n52556), .C0(n47341), .Z(n52557));
    PFUMX i40962 (.BLUT(n52552), .ALUT(n52553), .C0(n47341), .Z(n52554));
    PFUMX i40960 (.BLUT(n52549), .ALUT(n52550), .C0(n47341), .Z(n52551));
    PFUMX i40958 (.BLUT(n52546), .ALUT(n52547), .C0(n47341), .Z(n52548));
    PFUMX i40956 (.BLUT(n52543), .ALUT(n52544), .C0(n47341), .Z(n52545));
    FD1P3IX tx_cnt_i2 (.D(tx_cnt_2__N_5022[2]), .SP(sys_clk_enable_238), 
            .CD(n52186), .CK(sys_clk), .Q(tx_cnt[2])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=7, LSE_RCOL=4, LSE_LLINE=283, LSE_RLINE=300 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam tx_cnt_i2.GSR = "ENABLED";
    FD1P3IX tx_cnt_i1 (.D(tx_cnt_2__N_5022[1]), .SP(sys_clk_enable_238), 
            .CD(n52186), .CK(sys_clk), .Q(tx_cnt[1])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=7, LSE_RCOL=4, LSE_LLINE=283, LSE_RLINE=300 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam tx_cnt_i1.GSR = "ENABLED";
    FD1P3AX tx_state_i2 (.D(tx_state_2__N_4950[2]), .SP(sys_clk_enable_239), 
            .CK(sys_clk), .Q(tx_state[2])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=7, LSE_RCOL=4, LSE_LLINE=283, LSE_RLINE=300 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam tx_state_i2.GSR = "ENABLED";
    FD1P3AX tx_state_i1 (.D(tx_state_2__N_4950[1]), .SP(sys_clk_enable_239), 
            .CK(sys_clk), .Q(tx_state[1])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=7, LSE_RCOL=4, LSE_LLINE=283, LSE_RLINE=300 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam tx_state_i1.GSR = "ENABLED";
    FD1P3IX counter_i0_i15 (.D(n1[15]), .SP(sys_clk_enable_237), .CD(n30763), 
            .CK(sys_clk), .Q(counter[15])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=7, LSE_RCOL=4, LSE_LLINE=283, LSE_RLINE=300 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam counter_i0_i15.GSR = "ENABLED";
    FD1P3IX counter_i0_i14 (.D(n1[14]), .SP(sys_clk_enable_237), .CD(n30763), 
            .CK(sys_clk), .Q(counter[14])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=7, LSE_RCOL=4, LSE_LLINE=283, LSE_RLINE=300 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam counter_i0_i14.GSR = "ENABLED";
    FD1P3IX counter_i0_i13 (.D(n1[13]), .SP(sys_clk_enable_237), .CD(n30763), 
            .CK(sys_clk), .Q(counter[13])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=7, LSE_RCOL=4, LSE_LLINE=283, LSE_RLINE=300 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam counter_i0_i13.GSR = "ENABLED";
    FD1P3IX counter_i0_i12 (.D(n1[12]), .SP(sys_clk_enable_237), .CD(n30763), 
            .CK(sys_clk), .Q(counter[12])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=7, LSE_RCOL=4, LSE_LLINE=283, LSE_RLINE=300 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam counter_i0_i12.GSR = "ENABLED";
    FD1P3IX counter_i0_i11 (.D(n1[11]), .SP(sys_clk_enable_237), .CD(n30763), 
            .CK(sys_clk), .Q(counter[11])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=7, LSE_RCOL=4, LSE_LLINE=283, LSE_RLINE=300 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam counter_i0_i11.GSR = "ENABLED";
    FD1P3IX counter_i0_i10 (.D(n1[10]), .SP(sys_clk_enable_237), .CD(n30763), 
            .CK(sys_clk), .Q(counter[10])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=7, LSE_RCOL=4, LSE_LLINE=283, LSE_RLINE=300 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam counter_i0_i10.GSR = "ENABLED";
    FD1P3IX counter_i0_i9 (.D(n1[9]), .SP(sys_clk_enable_237), .CD(n30763), 
            .CK(sys_clk), .Q(counter[9])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=7, LSE_RCOL=4, LSE_LLINE=283, LSE_RLINE=300 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam counter_i0_i9.GSR = "ENABLED";
    FD1P3AY tx_output_128 (.D(tx_output_N_5048), .SP(sys_clk_enable_237), 
            .CK(sys_clk), .Q(tx_output)) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=7, LSE_RCOL=4, LSE_LLINE=283, LSE_RLINE=300 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam tx_output_128.GSR = "ENABLED";
    FD1P3IX tx_cnt_i0 (.D(tx_cnt_2__N_5022[0]), .SP(sys_clk_enable_238), 
            .CD(n52186), .CK(sys_clk), .Q(tx_cnt[0])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=7, LSE_RCOL=4, LSE_LLINE=283, LSE_RLINE=300 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam tx_cnt_i0.GSR = "ENABLED";
    FD1P3AX tx_state_i0 (.D(tx_state_2__N_4950[0]), .SP(sys_clk_enable_239), 
            .CK(sys_clk), .Q(tx_state[0])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=7, LSE_RCOL=4, LSE_LLINE=283, LSE_RLINE=300 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/txmitt.v(286[11] 393[9])
    defparam tx_state_i0.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module \rxcver(FIFO=0) 
//

module \rxcver(FIFO=0)  (parity_en, sys_clk, sin_c, rx_rdy, rbr_rd, 
            n53885, databits, GND_net, \divisor[8] , \divisor[4] , 
            \divisor[6] , \divisor[3] , \divisor[1] , \divisor[2] , 
            \divisor[0] ) /* synthesis syn_module_defined=1 */ ;
    input parity_en;
    input sys_clk;
    input sin_c;
    output rx_rdy;
    input rbr_rd;
    input n53885;
    input [1:0]databits;
    input GND_net;
    input \divisor[8] ;
    input \divisor[4] ;
    input \divisor[6] ;
    input \divisor[3] ;
    input \divisor[1] ;
    input \divisor[2] ;
    input \divisor[0] ;
    
    wire sys_clk /* synthesis SET_AS_NETWORK=sys_clk, is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(220[10:17])
    
    wire n3, n109;
    wire [2:0]cs_state;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(136[17:25])
    
    wire n52535, n52534, sin_d0, sin_d0_delay, rx_idle_d1, rx_idle, 
        rx_idle_N_4909, rbr_7__N_4884;
    wire [3:0]databit_recved_num;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(104[29:47])
    
    wire n50929, n52185;
    wire [3:0]databit_recved_num_3__N_4824;
    
    wire n43885;
    wire [15:0]counter;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(148[17:24])
    
    wire n15171;
    wire [15:0]n69;
    
    wire n43884, n43883, n43882, n43881;
    wire [15:0]n86;
    
    wire n43880, n43879, n43878, n47049, n39524, n49514, sys_clk_enable_240;
    wire [2:0]cs_state_2__N_4770;
    
    wire hunt_one_N_4910, n23, n21, n10, sys_clk_enable_156, n6715, 
        n30801, n43719, n43720, n34217, sys_clk_enable_241, n39528, 
        sys_clk_enable_171;
    wire [15:0]n87;
    
    wire n17, n30_adj_5095, n26_adj_5096, n18, n28_adj_5097, n22, 
        n49271, n43721, n49371, n49373, n26_adj_5098, n49367, n49336, 
        n52536;
    
    LUT4 cs_state_0__bdd_3_lut_40860_4_lut_4_lut_then_4_lut (.A(n3), .B(n109), 
         .C(cs_state[0]), .D(cs_state[1]), .Z(n52535)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(136[17:25])
    defparam cs_state_0__bdd_3_lut_40860_4_lut_4_lut_then_4_lut.init = 16'h0008;
    LUT4 cs_state_0__bdd_3_lut_40860_4_lut_4_lut_else_4_lut (.A(parity_en), 
         .B(cs_state[0]), .C(cs_state[1]), .Z(n52534)) /* synthesis lut_function=(!(A (B+!(C))+!A (B (C)+!B !(C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(136[17:25])
    defparam cs_state_0__bdd_3_lut_40860_4_lut_4_lut_else_4_lut.init = 16'h3434;
    FD1S3AX sin_d0_165 (.D(sin_c), .CK(sys_clk), .Q(sin_d0)) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=6, LSE_RCOL=4, LSE_LLINE=259, LSE_RLINE=279 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(455[14] 461[14])
    defparam sin_d0_165.GSR = "ENABLED";
    FD1S3AX sin_d0_delay_166 (.D(sin_d0), .CK(sys_clk), .Q(sin_d0_delay)) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=6, LSE_RCOL=4, LSE_LLINE=259, LSE_RLINE=279 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(455[14] 461[14])
    defparam sin_d0_delay_166.GSR = "ENABLED";
    FD1S3AY rx_idle_d1_169 (.D(rx_idle), .CK(sys_clk), .Q(rx_idle_d1)) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=6, LSE_RCOL=4, LSE_LLINE=259, LSE_RLINE=279 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(483[14] 486[14])
    defparam rx_idle_d1_169.GSR = "ENABLED";
    FD1S3AY rx_idle_157 (.D(rx_idle_N_4909), .CK(sys_clk), .Q(rx_idle)) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=6, LSE_RCOL=4, LSE_LLINE=259, LSE_RLINE=279 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(252[11] 255[27])
    defparam rx_idle_157.GSR = "ENABLED";
    FD1P3IX rbr_datardy_154 (.D(n53885), .SP(rbr_7__N_4884), .CD(rbr_rd), 
            .CK(sys_clk), .Q(rx_rdy)) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=6, LSE_RCOL=4, LSE_LLINE=259, LSE_RLINE=279 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(219[14] 227[12])
    defparam rbr_datardy_154.GSR = "ENABLED";
    LUT4 databits_0__bdd_4_lut_40566 (.A(databits[0]), .B(databit_recved_num[1]), 
         .C(databit_recved_num[0]), .D(databits[1]), .Z(n50929)) /* synthesis lut_function=(!(A ((C+(D))+!B)+!A !(B (C (D))+!B !((D)+!C)))) */ ;
    defparam databits_0__bdd_4_lut_40566.init = 16'h4018;
    LUT4 i25_3_lut_4_lut (.A(databit_recved_num[1]), .B(n52185), .C(databit_recved_num[3]), 
         .D(databit_recved_num[2]), .Z(databit_recved_num_3__N_4824[3])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(326[45:70])
    defparam i25_3_lut_4_lut.init = 16'h78f0;
    CCU2D counter_6620_add_4_17 (.A0(counter[15]), .B0(n15171), .C0(GND_net), 
          .D0(GND_net), .A1(GND_net), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n43885), .S0(n69[15]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620_add_4_17.INIT0 = 16'h7777;
    defparam counter_6620_add_4_17.INIT1 = 16'h0000;
    defparam counter_6620_add_4_17.INJECT1_0 = "NO";
    defparam counter_6620_add_4_17.INJECT1_1 = "NO";
    CCU2D counter_6620_add_4_15 (.A0(counter[13]), .B0(n15171), .C0(GND_net), 
          .D0(GND_net), .A1(counter[14]), .B1(n15171), .C1(GND_net), 
          .D1(GND_net), .CIN(n43884), .COUT(n43885), .S0(n69[13]), .S1(n69[14]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620_add_4_15.INIT0 = 16'h7777;
    defparam counter_6620_add_4_15.INIT1 = 16'h7777;
    defparam counter_6620_add_4_15.INJECT1_0 = "NO";
    defparam counter_6620_add_4_15.INJECT1_1 = "NO";
    CCU2D counter_6620_add_4_13 (.A0(counter[11]), .B0(n15171), .C0(GND_net), 
          .D0(GND_net), .A1(counter[12]), .B1(n15171), .C1(GND_net), 
          .D1(GND_net), .CIN(n43883), .COUT(n43884), .S0(n69[11]), .S1(n69[12]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620_add_4_13.INIT0 = 16'h7777;
    defparam counter_6620_add_4_13.INIT1 = 16'h7777;
    defparam counter_6620_add_4_13.INJECT1_0 = "NO";
    defparam counter_6620_add_4_13.INJECT1_1 = "NO";
    CCU2D counter_6620_add_4_11 (.A0(counter[9]), .B0(n15171), .C0(GND_net), 
          .D0(GND_net), .A1(counter[10]), .B1(n15171), .C1(GND_net), 
          .D1(GND_net), .CIN(n43882), .COUT(n43883), .S0(n69[9]), .S1(n69[10]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620_add_4_11.INIT0 = 16'h7777;
    defparam counter_6620_add_4_11.INIT1 = 16'h7777;
    defparam counter_6620_add_4_11.INJECT1_0 = "NO";
    defparam counter_6620_add_4_11.INJECT1_1 = "NO";
    CCU2D counter_6620_add_4_9 (.A0(counter[7]), .B0(n15171), .C0(GND_net), 
          .D0(GND_net), .A1(n86[8]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n43881), .COUT(n43882), .S0(n69[7]), .S1(n69[8]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620_add_4_9.INIT0 = 16'h7777;
    defparam counter_6620_add_4_9.INIT1 = 16'h0555;
    defparam counter_6620_add_4_9.INJECT1_0 = "NO";
    defparam counter_6620_add_4_9.INJECT1_1 = "NO";
    CCU2D counter_6620_add_4_7 (.A0(n86[5]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n86[6]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n43880), .COUT(n43881), .S0(n69[5]), .S1(n69[6]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620_add_4_7.INIT0 = 16'h0555;
    defparam counter_6620_add_4_7.INIT1 = 16'h0555;
    defparam counter_6620_add_4_7.INJECT1_0 = "NO";
    defparam counter_6620_add_4_7.INJECT1_1 = "NO";
    CCU2D counter_6620_add_4_5 (.A0(n86[3]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n86[4]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n43879), .COUT(n43880), .S0(n69[3]), .S1(n69[4]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620_add_4_5.INIT0 = 16'h0555;
    defparam counter_6620_add_4_5.INIT1 = 16'h0555;
    defparam counter_6620_add_4_5.INJECT1_0 = "NO";
    defparam counter_6620_add_4_5.INJECT1_1 = "NO";
    CCU2D counter_6620_add_4_3 (.A0(n86[1]), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n86[2]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .CIN(n43878), .COUT(n43879), .S0(n69[1]), .S1(n69[2]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620_add_4_3.INIT0 = 16'h0555;
    defparam counter_6620_add_4_3.INIT1 = 16'h0555;
    defparam counter_6620_add_4_3.INJECT1_0 = "NO";
    defparam counter_6620_add_4_3.INJECT1_1 = "NO";
    CCU2D counter_6620_add_4_1 (.A0(GND_net), .B0(GND_net), .C0(GND_net), 
          .D0(GND_net), .A1(n86[0]), .B1(GND_net), .C1(GND_net), .D1(GND_net), 
          .COUT(n43878), .S1(n69[0]));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620_add_4_1.INIT0 = 16'hF000;
    defparam counter_6620_add_4_1.INIT1 = 16'h0555;
    defparam counter_6620_add_4_1.INJECT1_0 = "NO";
    defparam counter_6620_add_4_1.INJECT1_1 = "NO";
    LUT4 i24_4_lut_3_lut (.A(cs_state[2]), .B(cs_state[1]), .C(cs_state[0]), 
         .Z(n47049)) /* synthesis lut_function=(!(A (B+(C))+!A (B (C)+!B !(C)))) */ ;
    defparam i24_4_lut_3_lut.init = 16'h1616;
    LUT4 i1_4_lut (.A(cs_state[2]), .B(n39524), .C(n49514), .D(cs_state[0]), 
         .Z(sys_clk_enable_240)) /* synthesis lut_function=(A+(B (C+!(D))+!B (C (D)))) */ ;
    defparam i1_4_lut.init = 16'hfaee;
    LUT4 i26649_3_lut (.A(cs_state[0]), .B(cs_state[2]), .C(cs_state[1]), 
         .Z(cs_state_2__N_4770[1])) /* synthesis lut_function=(!(A (B+(C))+!A (B+!(C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam i26649_3_lut.init = 16'h1212;
    LUT4 i28906_4_lut (.A(sin_d0), .B(n3), .C(cs_state[1]), .D(sin_d0_delay), 
         .Z(n39524)) /* synthesis lut_function=(A (B (C))+!A (B (C+(D))+!B !(C+!(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(136[17:25])
    defparam i28906_4_lut.init = 16'hc5c0;
    LUT4 i38719_4_lut (.A(n3), .B(hunt_one_N_4910), .C(cs_state[1]), .D(n23), 
         .Z(n49514)) /* synthesis lut_function=(A (B (C+(D))+!B !(C+!(D)))+!A (B (C))) */ ;
    defparam i38719_4_lut.init = 16'hcac0;
    LUT4 i1_4_lut_adj_141 (.A(databit_recved_num[0]), .B(n21), .C(n10), 
         .D(databits[1]), .Z(n23)) /* synthesis lut_function=(A (B)+!A (B+!(C+!(D)))) */ ;
    defparam i1_4_lut_adj_141.init = 16'hcdcc;
    LUT4 i1_3_lut (.A(databit_recved_num[2]), .B(databit_recved_num[3]), 
         .C(n50929), .Z(n21)) /* synthesis lut_function=(!((B+!(C))+!A)) */ ;
    defparam i1_3_lut.init = 16'h2020;
    LUT4 i39899_2_lut_3_lut (.A(cs_state[0]), .B(cs_state[1]), .C(cs_state[2]), 
         .Z(rx_idle_N_4909)) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam i39899_2_lut_3_lut.init = 16'h0101;
    LUT4 i39716_2_lut_rep_315_3_lut (.A(cs_state[0]), .B(cs_state[1]), .C(cs_state[2]), 
         .Z(sys_clk_enable_156)) /* synthesis lut_function=(!(A (C)+!A (B (C)))) */ ;
    defparam i39716_2_lut_rep_315_3_lut.init = 16'h1f1f;
    LUT4 i20129_2_lut_3_lut_4_lut (.A(cs_state[0]), .B(cs_state[1]), .C(n6715), 
         .D(cs_state[2]), .Z(n30801)) /* synthesis lut_function=(!(A ((D)+!C)+!A (B ((D)+!C)+!B !(C)))) */ ;
    defparam i20129_2_lut_3_lut_4_lut.init = 16'h10f0;
    LUT4 i2_4_lut (.A(cs_state[1]), .B(hunt_one_N_4910), .C(n3), .D(sin_d0), 
         .Z(n109)) /* synthesis lut_function=(A+(B (C+(D))+!B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(136[17:25])
    defparam i2_4_lut.init = 16'hfefa;
    CCU2D counter_15__I_0_13 (.A0(counter[14]), .B0(counter[13]), .C0(counter[12]), 
          .D0(counter[11]), .A1(counter[10]), .B1(counter[9]), .C1(counter[8]), 
          .D1(counter[6]), .CIN(n43719), .COUT(n43720));
    defparam counter_15__I_0_13.INIT0 = 16'h0001;
    defparam counter_15__I_0_13.INIT1 = 16'h0001;
    defparam counter_15__I_0_13.INJECT1_0 = "YES";
    defparam counter_15__I_0_13.INJECT1_1 = "YES";
    LUT4 i1_3_lut_4_lut (.A(cs_state[2]), .B(cs_state[1]), .C(n34217), 
         .D(cs_state[0]), .Z(sys_clk_enable_241)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (C+(D)))) */ ;
    defparam i1_3_lut_4_lut.init = 16'hf1f0;
    LUT4 i28920_4_lut_4_lut (.A(cs_state[2]), .B(cs_state[0]), .C(n39528), 
         .D(n39524), .Z(sys_clk_enable_171)) /* synthesis lut_function=(A (C)+!A (B (C)+!B (D))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(136[17:25])
    defparam i28920_4_lut_4_lut.init = 16'hf1e0;
    LUT4 i7616_2_lut_3_lut_4_lut (.A(databit_recved_num[0]), .B(hunt_one_N_4910), 
         .C(databit_recved_num[2]), .D(databit_recved_num[1]), .Z(databit_recved_num_3__N_4824[2])) /* synthesis lut_function=(!(A (B (C (D)+!C !(D))+!B !(C))+!A !(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(326[45:70])
    defparam i7616_2_lut_3_lut_4_lut.init = 16'h78f0;
    LUT4 rx_idle_I_0_188_2_lut (.A(rx_idle), .B(rx_idle_d1), .Z(rbr_7__N_4884)) /* synthesis lut_function=(!((B)+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(437[18:59])
    defparam rx_idle_I_0_188_2_lut.init = 16'h2222;
    FD1P3AX counter_6620__i0 (.D(n87[0]), .SP(sys_clk_enable_156), .CK(sys_clk), 
            .Q(counter[0])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620__i0.GSR = "ENABLED";
    LUT4 i28953_4_lut (.A(n3), .B(cs_state[2]), .C(cs_state[0]), .D(cs_state[1]), 
         .Z(n15171)) /* synthesis lut_function=(!(A (B+!(C (D)))+!A (B (C+(D))+!B !(C+(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(136[17:25])
    defparam i28953_4_lut.init = 16'h3114;
    LUT4 i39870_4_lut (.A(n17), .B(n30_adj_5095), .C(n26_adj_5096), .D(n18), 
         .Z(n3)) /* synthesis lut_function=(!(A+(B+(C+(D))))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(136[17:25])
    defparam i39870_4_lut.init = 16'h0001;
    LUT4 i1_2_lut (.A(counter[0]), .B(counter[14]), .Z(n17)) /* synthesis lut_function=((B)+!A) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(313[20:54])
    defparam i1_2_lut.init = 16'hdddd;
    LUT4 i14_4_lut (.A(counter[2]), .B(n28_adj_5097), .C(n22), .D(counter[4]), 
         .Z(n30_adj_5095)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(313[20:54])
    defparam i14_4_lut.init = 16'hfffe;
    LUT4 i10_4_lut (.A(counter[8]), .B(counter[7]), .C(counter[10]), .D(counter[1]), 
         .Z(n26_adj_5096)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(313[20:54])
    defparam i10_4_lut.init = 16'hfffe;
    LUT4 i2_2_lut (.A(counter[9]), .B(counter[3]), .Z(n18)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(313[20:54])
    defparam i2_2_lut.init = 16'heeee;
    LUT4 i12_4_lut (.A(counter[11]), .B(counter[13]), .C(counter[5]), 
         .D(counter[6]), .Z(n28_adj_5097)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(313[20:54])
    defparam i12_4_lut.init = 16'hfffe;
    LUT4 i6_2_lut (.A(counter[12]), .B(counter[15]), .Z(n22)) /* synthesis lut_function=(A+(B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(313[20:54])
    defparam i6_2_lut.init = 16'heeee;
    LUT4 counter_6620_mux_5_i9_3_lut (.A(\divisor[8] ), .B(counter[8]), 
         .C(n15171), .Z(n86[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620_mux_5_i9_3_lut.init = 16'hcaca;
    LUT4 counter_6620_mux_5_i6_3_lut (.A(\divisor[4] ), .B(counter[5]), 
         .C(n15171), .Z(n86[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620_mux_5_i6_3_lut.init = 16'hcaca;
    LUT4 counter_6620_mux_5_i7_3_lut (.A(\divisor[6] ), .B(counter[6]), 
         .C(n15171), .Z(n86[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620_mux_5_i7_3_lut.init = 16'hcaca;
    LUT4 counter_6620_mux_5_i4_3_lut (.A(\divisor[3] ), .B(counter[3]), 
         .C(n15171), .Z(n86[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620_mux_5_i4_3_lut.init = 16'hcaca;
    LUT4 counter_6620_mux_5_i5_3_lut (.A(\divisor[4] ), .B(counter[4]), 
         .C(n15171), .Z(n86[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620_mux_5_i5_3_lut.init = 16'hcaca;
    LUT4 counter_6620_mux_5_i2_3_lut (.A(\divisor[1] ), .B(counter[1]), 
         .C(n15171), .Z(n86[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620_mux_5_i2_3_lut.init = 16'hcaca;
    LUT4 counter_6620_mux_5_i3_3_lut (.A(\divisor[2] ), .B(counter[2]), 
         .C(n15171), .Z(n86[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620_mux_5_i3_3_lut.init = 16'hcaca;
    LUT4 counter_6620_mux_6_i2_3_lut (.A(n69[1]), .B(\divisor[1] ), .C(n6715), 
         .Z(n87[1])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620_mux_6_i2_3_lut.init = 16'hcaca;
    LUT4 counter_6620_mux_6_i3_3_lut (.A(n69[2]), .B(\divisor[2] ), .C(n6715), 
         .Z(n87[2])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620_mux_6_i3_3_lut.init = 16'hcaca;
    LUT4 counter_6620_mux_6_i4_3_lut (.A(n69[3]), .B(\divisor[3] ), .C(n6715), 
         .Z(n87[3])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620_mux_6_i4_3_lut.init = 16'hcaca;
    LUT4 counter_6620_mux_6_i5_3_lut (.A(n69[4]), .B(\divisor[4] ), .C(n6715), 
         .Z(n87[4])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620_mux_6_i5_3_lut.init = 16'hcaca;
    LUT4 counter_6620_mux_6_i6_3_lut (.A(n69[5]), .B(\divisor[4] ), .C(n6715), 
         .Z(n87[5])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620_mux_6_i6_3_lut.init = 16'hcaca;
    LUT4 counter_6620_mux_6_i7_3_lut (.A(n69[6]), .B(\divisor[6] ), .C(n6715), 
         .Z(n87[6])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620_mux_6_i7_3_lut.init = 16'hcaca;
    LUT4 counter_6620_mux_6_i9_3_lut (.A(n69[8]), .B(\divisor[8] ), .C(n6715), 
         .Z(n87[8])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620_mux_6_i9_3_lut.init = 16'hcaca;
    LUT4 i28910_4_lut (.A(n109), .B(cs_state[2]), .C(cs_state[0]), .D(n49514), 
         .Z(n39528)) /* synthesis lut_function=(A (B+((D)+!C))+!A (B (C)+!B (C (D)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(136[17:25])
    defparam i28910_4_lut.init = 16'hfaca;
    LUT4 i39946_3_lut (.A(cs_state[1]), .B(cs_state[2]), .C(cs_state[0]), 
         .Z(cs_state_2__N_4770[2])) /* synthesis lut_function=(!(A+(B+(C)))) */ ;
    defparam i39946_3_lut.init = 16'h0101;
    LUT4 i4_4_lut (.A(hunt_one_N_4910), .B(cs_state[1]), .C(cs_state[2]), 
         .D(n49271), .Z(n34217)) /* synthesis lut_function=(!((B+((D)+!C))+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(136[17:25])
    defparam i4_4_lut.init = 16'h0020;
    LUT4 i38479_2_lut (.A(cs_state[0]), .B(sin_d0), .Z(n49271)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i38479_2_lut.init = 16'heeee;
    LUT4 counter_6620_mux_5_i1_3_lut (.A(\divisor[0] ), .B(counter[0]), 
         .C(n15171), .Z(n86[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620_mux_5_i1_3_lut.init = 16'hcaca;
    LUT4 i7603_2_lut_rep_249 (.A(databit_recved_num[0]), .B(hunt_one_N_4910), 
         .Z(n52185)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(326[45:70])
    defparam i7603_2_lut_rep_249.init = 16'h8888;
    FD1P3AX cs_state_i1 (.D(cs_state_2__N_4770[1]), .SP(sys_clk_enable_240), 
            .CK(sys_clk), .Q(cs_state[1])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=6, LSE_RCOL=4, LSE_LLINE=259, LSE_RLINE=279 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam cs_state_i1.GSR = "ENABLED";
    LUT4 i7601_2_lut (.A(databit_recved_num[0]), .B(hunt_one_N_4910), .Z(databit_recved_num_3__N_4824[0])) /* synthesis lut_function=(!(A (B)+!A !(B))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(326[45:70])
    defparam i7601_2_lut.init = 16'h6666;
    CCU2D counter_15__I_0_0 (.A0(\divisor[8] ), .B0(counter[7]), .C0(GND_net), 
          .D0(GND_net), .A1(counter[15]), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .COUT(n43719));   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(186[39:61])
    defparam counter_15__I_0_0.INIT0 = 16'h9000;
    defparam counter_15__I_0_0.INIT1 = 16'h5555;
    defparam counter_15__I_0_0.INJECT1_0 = "NO";
    defparam counter_15__I_0_0.INJECT1_1 = "YES";
    LUT4 i7609_2_lut_3_lut (.A(databit_recved_num[0]), .B(hunt_one_N_4910), 
         .C(databit_recved_num[1]), .Z(databit_recved_num_3__N_4824[1])) /* synthesis lut_function=(!(A (B (C)+!B !(C))+!A !(C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(326[45:70])
    defparam i7609_2_lut_3_lut.init = 16'h7878;
    CCU2D counter_15__I_0_16 (.A0(\divisor[2] ), .B0(counter[1]), .C0(\divisor[1] ), 
          .D0(counter[0]), .A1(GND_net), .B1(GND_net), .C1(GND_net), 
          .D1(GND_net), .CIN(n43721), .S1(hunt_one_N_4910));
    defparam counter_15__I_0_16.INIT0 = 16'h9009;
    defparam counter_15__I_0_16.INIT1 = 16'hFFFF;
    defparam counter_15__I_0_16.INJECT1_0 = "YES";
    defparam counter_15__I_0_16.INJECT1_1 = "NO";
    LUT4 i4_4_lut_4_lut (.A(databits[0]), .B(databit_recved_num[1]), .C(databit_recved_num[2]), 
         .D(databit_recved_num[3]), .Z(n10)) /* synthesis lut_function=((B+(C+!(D)))+!A) */ ;
    defparam i4_4_lut_4_lut.init = 16'hfdff;
    LUT4 counter_6620_mux_6_i1_3_lut (.A(n69[0]), .B(\divisor[0] ), .C(n6715), 
         .Z(n87[0])) /* synthesis lut_function=(A (B+!(C))+!A (B (C))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620_mux_6_i1_3_lut.init = 16'hcaca;
    LUT4 i1_4_lut_adj_142 (.A(counter[0]), .B(n49371), .C(n49373), .D(n26_adj_5098), 
         .Z(n6715)) /* synthesis lut_function=(!((B+(C+!(D)))+!A)) */ ;
    defparam i1_4_lut_adj_142.init = 16'h0200;
    LUT4 i38576_4_lut (.A(counter[9]), .B(counter[5]), .C(counter[8]), 
         .D(counter[13]), .Z(n49371)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i38576_4_lut.init = 16'hfffe;
    LUT4 i38578_4_lut (.A(counter[7]), .B(n49367), .C(n49336), .D(counter[10]), 
         .Z(n49373)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i38578_4_lut.init = 16'hfffe;
    LUT4 i10_4_lut_adj_143 (.A(n47049), .B(counter[3]), .C(counter[2]), 
         .D(counter[6]), .Z(n26_adj_5098)) /* synthesis lut_function=(!((B+(C+(D)))+!A)) */ ;
    defparam i10_4_lut_adj_143.init = 16'h0002;
    LUT4 i38572_4_lut (.A(counter[12]), .B(counter[4]), .C(counter[1]), 
         .D(counter[14]), .Z(n49367)) /* synthesis lut_function=(A+(B+(C+(D)))) */ ;
    defparam i38572_4_lut.init = 16'hfffe;
    LUT4 i38541_2_lut (.A(counter[15]), .B(counter[11]), .Z(n49336)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i38541_2_lut.init = 16'heeee;
    FD1P3AX counter_6620__i1 (.D(n87[1]), .SP(sys_clk_enable_156), .CK(sys_clk), 
            .Q(counter[1])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620__i1.GSR = "ENABLED";
    FD1P3AX counter_6620__i2 (.D(n87[2]), .SP(sys_clk_enable_156), .CK(sys_clk), 
            .Q(counter[2])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620__i2.GSR = "ENABLED";
    FD1P3AX counter_6620__i3 (.D(n87[3]), .SP(sys_clk_enable_156), .CK(sys_clk), 
            .Q(counter[3])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620__i3.GSR = "ENABLED";
    FD1P3AX counter_6620__i4 (.D(n87[4]), .SP(sys_clk_enable_156), .CK(sys_clk), 
            .Q(counter[4])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620__i4.GSR = "ENABLED";
    FD1P3AX counter_6620__i5 (.D(n87[5]), .SP(sys_clk_enable_156), .CK(sys_clk), 
            .Q(counter[5])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620__i5.GSR = "ENABLED";
    FD1P3AX counter_6620__i6 (.D(n87[6]), .SP(sys_clk_enable_156), .CK(sys_clk), 
            .Q(counter[6])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620__i6.GSR = "ENABLED";
    FD1P3AX counter_6620__i8 (.D(n87[8]), .SP(sys_clk_enable_156), .CK(sys_clk), 
            .Q(counter[8])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620__i8.GSR = "ENABLED";
    CCU2D counter_15__I_0_15 (.A0(\divisor[6] ), .B0(counter[5]), .C0(\divisor[4] ), 
          .D0(counter[4]), .A1(\divisor[4] ), .B1(counter[3]), .C1(\divisor[3] ), 
          .D1(counter[2]), .CIN(n43720), .COUT(n43721));
    defparam counter_15__I_0_15.INIT0 = 16'h9009;
    defparam counter_15__I_0_15.INIT1 = 16'h9009;
    defparam counter_15__I_0_15.INJECT1_0 = "YES";
    defparam counter_15__I_0_15.INJECT1_1 = "YES";
    PFUMX i40950 (.BLUT(n52534), .ALUT(n52535), .C0(cs_state[2]), .Z(n52536));
    FD1P3IX counter_6620__i15 (.D(n69[15]), .SP(sys_clk_enable_156), .CD(n30801), 
            .CK(sys_clk), .Q(counter[15])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620__i15.GSR = "ENABLED";
    FD1P3IX counter_6620__i14 (.D(n69[14]), .SP(sys_clk_enable_156), .CD(n30801), 
            .CK(sys_clk), .Q(counter[14])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620__i14.GSR = "ENABLED";
    FD1P3IX counter_6620__i13 (.D(n69[13]), .SP(sys_clk_enable_156), .CD(n30801), 
            .CK(sys_clk), .Q(counter[13])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620__i13.GSR = "ENABLED";
    FD1P3IX counter_6620__i12 (.D(n69[12]), .SP(sys_clk_enable_156), .CD(n30801), 
            .CK(sys_clk), .Q(counter[12])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620__i12.GSR = "ENABLED";
    FD1P3IX counter_6620__i11 (.D(n69[11]), .SP(sys_clk_enable_156), .CD(n30801), 
            .CK(sys_clk), .Q(counter[11])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620__i11.GSR = "ENABLED";
    FD1P3IX counter_6620__i10 (.D(n69[10]), .SP(sys_clk_enable_156), .CD(n30801), 
            .CK(sys_clk), .Q(counter[10])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620__i10.GSR = "ENABLED";
    FD1P3IX counter_6620__i9 (.D(n69[9]), .SP(sys_clk_enable_156), .CD(n30801), 
            .CK(sys_clk), .Q(counter[9])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620__i9.GSR = "ENABLED";
    FD1P3IX counter_6620__i7 (.D(n69[7]), .SP(sys_clk_enable_156), .CD(n30801), 
            .CK(sys_clk), .Q(counter[7])) /* synthesis syn_use_carry_chain=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam counter_6620__i7.GSR = "ENABLED";
    FD1P3AX cs_state_i2 (.D(cs_state_2__N_4770[2]), .SP(sys_clk_enable_171), 
            .CK(sys_clk), .Q(cs_state[2])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=6, LSE_RCOL=4, LSE_LLINE=259, LSE_RLINE=279 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam cs_state_i2.GSR = "ENABLED";
    FD1P3IX databit_recved_num_i3 (.D(databit_recved_num_3__N_4824[3]), .SP(sys_clk_enable_241), 
            .CD(n34217), .CK(sys_clk), .Q(databit_recved_num[3])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=6, LSE_RCOL=4, LSE_LLINE=259, LSE_RLINE=279 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam databit_recved_num_i3.GSR = "ENABLED";
    FD1P3IX databit_recved_num_i2 (.D(databit_recved_num_3__N_4824[2]), .SP(sys_clk_enable_241), 
            .CD(n34217), .CK(sys_clk), .Q(databit_recved_num[2])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=6, LSE_RCOL=4, LSE_LLINE=259, LSE_RLINE=279 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam databit_recved_num_i2.GSR = "ENABLED";
    FD1P3IX databit_recved_num_i1 (.D(databit_recved_num_3__N_4824[1]), .SP(sys_clk_enable_241), 
            .CD(n34217), .CK(sys_clk), .Q(databit_recved_num[1])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=6, LSE_RCOL=4, LSE_LLINE=259, LSE_RLINE=279 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam databit_recved_num_i1.GSR = "ENABLED";
    FD1P3AX cs_state_i0 (.D(n52536), .SP(sys_clk_enable_240), .CK(sys_clk), 
            .Q(cs_state[0])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=6, LSE_RCOL=4, LSE_LLINE=259, LSE_RLINE=279 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam cs_state_i0.GSR = "ENABLED";
    FD1P3IX databit_recved_num_i0 (.D(databit_recved_num_3__N_4824[0]), .SP(sys_clk_enable_241), 
            .CD(n34217), .CK(sys_clk), .Q(databit_recved_num[0])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=6, LSE_RCOL=4, LSE_LLINE=259, LSE_RLINE=279 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/rxcver.v(289[8] 376[18])
    defparam databit_recved_num_i0.GSR = "ENABLED";
    
endmodule
//
// Verilog Description of module \intface(CLK_IN_MHZ=38) 
//

module \intface(CLK_IN_MHZ=38)  (\adr_i[0] , cyc_i, we_i, \adr_i[1] , 
            \adr_i[2] , \THR[0] , sys_clk, \dat_i[0] , databits, \divisor[0] , 
            thr_wr, rbr_rd, \next_state_9__N_4541[6] , n53885, rx_rdy, 
            rxrdy_n_c, \THR[1] , \dat_i[1] , \THR[2] , \dat_i[2] , 
            \THR[3] , \dat_i[3] , \THR[4] , \dat_i[5] , \THR[6] , 
            \dat_i[6] , \lcr[2] , parity_en, parity_even, tx_break, 
            \divisor[1] , \divisor[2] , \divisor[3] , \divisor[4] , 
            \divisor[6] , \divisor[8] , n53884) /* synthesis syn_module_defined=1 */ ;
    input \adr_i[0] ;
    input cyc_i;
    input we_i;
    input \adr_i[1] ;
    input \adr_i[2] ;
    output \THR[0] ;
    input sys_clk;
    input \dat_i[0] ;
    output [1:0]databits;
    output \divisor[0] ;
    output thr_wr;
    output rbr_rd;
    output \next_state_9__N_4541[6] ;
    input n53885;
    input rx_rdy;
    output rxrdy_n_c;
    output \THR[1] ;
    input \dat_i[1] ;
    output \THR[2] ;
    input \dat_i[2] ;
    output \THR[3] ;
    input \dat_i[3] ;
    output \THR[4] ;
    input \dat_i[5] ;
    output \THR[6] ;
    input \dat_i[6] ;
    output \lcr[2] ;
    output parity_en;
    output parity_even;
    output tx_break;
    output \divisor[1] ;
    output \divisor[2] ;
    output \divisor[3] ;
    output \divisor[4] ;
    output \divisor[6] ;
    output \divisor[8] ;
    input n53884;
    
    wire sys_clk /* synthesis SET_AS_NETWORK=sys_clk, is_clock=1 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/drone2.v(220[10:17])
    
    wire n52397, rbr_rd_strobe, n52396, sys_clk_enable_140, div_wr_strobe, 
        sys_clk_enable_129, thr_wr_strobe;
    
    LUT4 i2_3_lut_4_lut (.A(\adr_i[0] ), .B(n52397), .C(cyc_i), .D(we_i), 
         .Z(rbr_rd_strobe)) /* synthesis lut_function=(!(A+(B+((D)+!C)))) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/intface.v(338[8:13])
    defparam i2_3_lut_4_lut.init = 16'h0010;
    LUT4 i1_2_lut_4_lut (.A(\adr_i[1] ), .B(n52396), .C(\adr_i[0] ), .D(\adr_i[2] ), 
         .Z(sys_clk_enable_140)) /* synthesis lut_function=(!((((D)+!C)+!B)+!A)) */ ;
    defparam i1_2_lut_4_lut.init = 16'h0080;
    LUT4 i1_2_lut_4_lut_adj_140 (.A(\adr_i[1] ), .B(n52396), .C(\adr_i[0] ), 
         .D(\adr_i[2] ), .Z(div_wr_strobe)) /* synthesis lut_function=(A (B (C (D)))) */ ;
    defparam i1_2_lut_4_lut_adj_140.init = 16'h8000;
    FD1P3AX thr_nonfifo_i0_i0 (.D(\dat_i[0] ), .SP(sys_clk_enable_129), 
            .CK(sys_clk), .Q(\THR[0] )) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=10, LSE_RCOL=4, LSE_LLINE=169, LSE_RLINE=209 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/intface.v(365[13] 376[18])
    defparam thr_nonfifo_i0_i0.GSR = "ENABLED";
    FD1P3AX lcr__i1 (.D(\dat_i[0] ), .SP(sys_clk_enable_140), .CK(sys_clk), 
            .Q(databits[0])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=10, LSE_RCOL=4, LSE_LLINE=169, LSE_RLINE=209 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/intface.v(365[13] 376[18])
    defparam lcr__i1.GSR = "ENABLED";
    FD1P3AY divisor_i0_i0 (.D(\dat_i[0] ), .SP(div_wr_strobe), .CK(sys_clk), 
            .Q(\divisor[0] )) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=10, LSE_RCOL=4, LSE_LLINE=169, LSE_RLINE=209 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/intface.v(230[12] 231[32])
    defparam divisor_i0_i0.GSR = "ENABLED";
    FD1S3AX thr_wr_138 (.D(thr_wr_strobe), .CK(sys_clk), .Q(thr_wr)) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=10, LSE_RCOL=4, LSE_LLINE=169, LSE_RLINE=209 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/intface.v(252[7:31])
    defparam thr_wr_138.GSR = "ENABLED";
    FD1S3AX rbr_rd_nonfifo_139 (.D(rbr_rd_strobe), .CK(sys_clk), .Q(rbr_rd)) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=10, LSE_RCOL=4, LSE_LLINE=169, LSE_RLINE=209 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/intface.v(263[6:38])
    defparam rbr_rd_nonfifo_139.GSR = "ENABLED";
    FD1P3IX ack_o_146 (.D(n53885), .SP(cyc_i), .CD(\next_state_9__N_4541[6] ), 
            .CK(sys_clk), .Q(\next_state_9__N_4541[6] )) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=10, LSE_RCOL=4, LSE_LLINE=169, LSE_RLINE=209 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/intface.v(629[10] 632[21])
    defparam ack_o_146.GSR = "ENABLED";
    LUT4 i1_2_lut_rep_460 (.A(cyc_i), .B(we_i), .Z(n52396)) /* synthesis lut_function=(A (B)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/intface.v(286[29:70])
    defparam i1_2_lut_rep_460.init = 16'h8888;
    LUT4 i3_3_lut_4_lut (.A(cyc_i), .B(we_i), .C(\adr_i[0] ), .D(n52397), 
         .Z(sys_clk_enable_129)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/intface.v(286[29:70])
    defparam i3_3_lut_4_lut.init = 16'h0008;
    LUT4 i1_2_lut_3_lut_4_lut (.A(cyc_i), .B(we_i), .C(n52397), .D(\adr_i[0] ), 
         .Z(thr_wr_strobe)) /* synthesis lut_function=(!(((C+(D))+!B)+!A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/intface.v(286[29:70])
    defparam i1_2_lut_3_lut_4_lut.init = 16'h0008;
    LUT4 i38554_2_lut_rep_461 (.A(\adr_i[1] ), .B(\adr_i[2] ), .Z(n52397)) /* synthesis lut_function=(A+(B)) */ ;
    defparam i38554_2_lut_rep_461.init = 16'heeee;
    LUT4 rx_rdy_I_0_1_lut (.A(rx_rdy), .Z(rxrdy_n_c)) /* synthesis lut_function=(!(A)) */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/uart_core.v(321[23:30])
    defparam rx_rdy_I_0_1_lut.init = 16'h5555;
    FD1P3AX thr_nonfifo_i0_i1 (.D(\dat_i[1] ), .SP(sys_clk_enable_129), 
            .CK(sys_clk), .Q(\THR[1] )) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=10, LSE_RCOL=4, LSE_LLINE=169, LSE_RLINE=209 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/intface.v(365[13] 376[18])
    defparam thr_nonfifo_i0_i1.GSR = "ENABLED";
    FD1P3AX thr_nonfifo_i0_i2 (.D(\dat_i[2] ), .SP(sys_clk_enable_129), 
            .CK(sys_clk), .Q(\THR[2] )) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=10, LSE_RCOL=4, LSE_LLINE=169, LSE_RLINE=209 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/intface.v(365[13] 376[18])
    defparam thr_nonfifo_i0_i2.GSR = "ENABLED";
    FD1P3AX thr_nonfifo_i0_i3 (.D(\dat_i[3] ), .SP(sys_clk_enable_129), 
            .CK(sys_clk), .Q(\THR[3] )) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=10, LSE_RCOL=4, LSE_LLINE=169, LSE_RLINE=209 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/intface.v(365[13] 376[18])
    defparam thr_nonfifo_i0_i3.GSR = "ENABLED";
    FD1P3AX thr_nonfifo_i0_i4 (.D(\dat_i[5] ), .SP(sys_clk_enable_129), 
            .CK(sys_clk), .Q(\THR[4] )) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=10, LSE_RCOL=4, LSE_LLINE=169, LSE_RLINE=209 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/intface.v(365[13] 376[18])
    defparam thr_nonfifo_i0_i4.GSR = "ENABLED";
    FD1P3AX thr_nonfifo_i0_i6 (.D(\dat_i[6] ), .SP(sys_clk_enable_129), 
            .CK(sys_clk), .Q(\THR[6] )) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=10, LSE_RCOL=4, LSE_LLINE=169, LSE_RLINE=209 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/intface.v(365[13] 376[18])
    defparam thr_nonfifo_i0_i6.GSR = "ENABLED";
    FD1P3AX lcr__i2 (.D(\dat_i[1] ), .SP(sys_clk_enable_140), .CK(sys_clk), 
            .Q(databits[1])) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=10, LSE_RCOL=4, LSE_LLINE=169, LSE_RLINE=209 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/intface.v(365[13] 376[18])
    defparam lcr__i2.GSR = "ENABLED";
    FD1P3AX lcr__i3 (.D(\dat_i[2] ), .SP(sys_clk_enable_140), .CK(sys_clk), 
            .Q(\lcr[2] )) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=10, LSE_RCOL=4, LSE_LLINE=169, LSE_RLINE=209 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/intface.v(365[13] 376[18])
    defparam lcr__i3.GSR = "ENABLED";
    FD1P3AX lcr__i4 (.D(\dat_i[3] ), .SP(sys_clk_enable_140), .CK(sys_clk), 
            .Q(parity_en)) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=10, LSE_RCOL=4, LSE_LLINE=169, LSE_RLINE=209 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/intface.v(365[13] 376[18])
    defparam lcr__i4.GSR = "ENABLED";
    FD1P3AX lcr__i5 (.D(\dat_i[5] ), .SP(sys_clk_enable_140), .CK(sys_clk), 
            .Q(parity_even)) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=10, LSE_RCOL=4, LSE_LLINE=169, LSE_RLINE=209 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/intface.v(365[13] 376[18])
    defparam lcr__i5.GSR = "ENABLED";
    FD1P3AX lcr__i7 (.D(\dat_i[6] ), .SP(sys_clk_enable_140), .CK(sys_clk), 
            .Q(tx_break)) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=10, LSE_RCOL=4, LSE_LLINE=169, LSE_RLINE=209 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/intface.v(365[13] 376[18])
    defparam lcr__i7.GSR = "ENABLED";
    FD1P3AX divisor_i0_i1 (.D(\dat_i[1] ), .SP(div_wr_strobe), .CK(sys_clk), 
            .Q(\divisor[1] )) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=10, LSE_RCOL=4, LSE_LLINE=169, LSE_RLINE=209 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/intface.v(230[12] 231[32])
    defparam divisor_i0_i1.GSR = "ENABLED";
    FD1P3AX divisor_i0_i2 (.D(\dat_i[2] ), .SP(div_wr_strobe), .CK(sys_clk), 
            .Q(\divisor[2] )) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=10, LSE_RCOL=4, LSE_LLINE=169, LSE_RLINE=209 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/intface.v(230[12] 231[32])
    defparam divisor_i0_i2.GSR = "ENABLED";
    FD1P3AY divisor_i0_i3 (.D(\dat_i[3] ), .SP(div_wr_strobe), .CK(sys_clk), 
            .Q(\divisor[3] )) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=10, LSE_RCOL=4, LSE_LLINE=169, LSE_RLINE=209 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/intface.v(230[12] 231[32])
    defparam divisor_i0_i3.GSR = "ENABLED";
    FD1P3AX divisor_i0_i4 (.D(\dat_i[5] ), .SP(div_wr_strobe), .CK(sys_clk), 
            .Q(\divisor[4] )) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=10, LSE_RCOL=4, LSE_LLINE=169, LSE_RLINE=209 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/intface.v(230[12] 231[32])
    defparam divisor_i0_i4.GSR = "ENABLED";
    FD1P3AY divisor_i0_i6 (.D(\dat_i[6] ), .SP(div_wr_strobe), .CK(sys_clk), 
            .Q(\divisor[6] )) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=10, LSE_RCOL=4, LSE_LLINE=169, LSE_RLINE=209 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/intface.v(230[12] 231[32])
    defparam divisor_i0_i6.GSR = "ENABLED";
    FD1P3AY divisor_i0_i8 (.D(n53884), .SP(div_wr_strobe), .CK(sys_clk), 
            .Q(\divisor[8] )) /* synthesis LSE_LINE_FILE_ID=24, LSE_LCOL=10, LSE_RCOL=4, LSE_LLINE=169, LSE_RLINE=209 */ ;   // c:/users/mintbox/documents/latticediamondprojects/ethans-fork-drone2-capstone/drone2_ls_capstone/source-code/drone2ethanfork/impl1/source/intface.v(230[12] 231[32])
    defparam divisor_i0_i8.GSR = "ENABLED";
    
endmodule
